* NGSPICE file created from basic.ext - technology: scmos

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

.subckt basic a gnd o vdd
X_2_ _1_/Y gnd o vdd BUFX2
X_1_ a gnd _1_/Y vdd INVX1
.ends

