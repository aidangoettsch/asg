* NGSPICE file created from mux_using_if.ext - technology: scmos

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

.subckt mux_using_if din_0 din_1 mux_out sel
X_5_ sel _5_/B _4_/Y _6_/gnd _6_/A _6_/vdd OAI21X1
X_6_ _6_/A _6_/gnd mux_out _6_/vdd BUFX2
X_3_ din_0 _6_/gnd _5_/B _6_/vdd INVX1
X_4_ din_1 sel _6_/gnd _4_/Y _6_/vdd NAND2X1
.ends

