VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO mux_using_if
   CLASS BLOCK ;
   FOREIGN mux_using_if ;
   ORIGIN 3.6000 -0.4000 ;
   SIZE 176.8000 BY 21.2000 ;
   PIN din_0
      PORT
         LAYER metal1 ;
	    RECT 18.8000 16.3000 19.6000 17.2000 ;
	    RECT 172.4000 16.3000 173.2000 16.4000 ;
	    RECT 18.8000 15.7000 173.2000 16.3000 ;
	    RECT 18.8000 15.6000 19.6000 15.7000 ;
	    RECT 172.4000 15.6000 173.2000 15.7000 ;
         LAYER metal2 ;
	    RECT 172.4000 17.6000 173.2000 18.4000 ;
	    RECT 172.5000 16.4000 173.1000 17.6000 ;
	    RECT 172.4000 15.6000 173.2000 16.4000 ;
         LAYER metal3 ;
	    RECT 172.4000 17.6000 173.2000 18.4000 ;
      END
   END din_0
   PIN din_1
      PORT
         LAYER metal1 ;
	    RECT 6.0000 13.6000 6.8000 15.2000 ;
         LAYER metal2 ;
	    RECT 6.0000 13.6000 6.8000 14.4000 ;
	    RECT 6.1000 10.4000 6.7000 13.6000 ;
	    RECT 6.0000 9.6000 6.8000 10.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 10.3000 6.8000 10.4000 ;
	    RECT -3.5000 9.7000 6.8000 10.3000 ;
	    RECT 6.0000 9.6000 6.8000 9.7000 ;
      END
   END din_1
   PIN mux_out
      PORT
         LAYER metal1 ;
	    RECT 1.2000 12.4000 2.0000 19.8000 ;
	    RECT 1.2000 10.2000 1.8000 12.4000 ;
	    RECT -3.6000 6.3000 -2.8000 6.4000 ;
	    RECT 1.2000 6.3000 2.0000 10.2000 ;
	    RECT -3.6000 5.7000 2.0000 6.3000 ;
	    RECT -3.6000 5.6000 -2.8000 5.7000 ;
	    RECT 1.2000 2.2000 2.0000 5.7000 ;
         LAYER metal2 ;
	    RECT -3.6000 5.6000 -2.8000 6.4000 ;
         LAYER metal3 ;
	    RECT -3.6000 5.6000 -2.8000 6.4000 ;
      END
   END mux_out
   PIN sel
      PORT
         LAYER metal1 ;
	    RECT 14.8000 14.4000 15.6000 14.8000 ;
	    RECT 14.8000 13.8000 16.4000 14.4000 ;
	    RECT 15.6000 13.6000 16.4000 13.8000 ;
	    RECT 9.2000 8.8000 10.0000 10.4000 ;
         LAYER metal2 ;
	    RECT 9.2000 13.6000 10.0000 14.4000 ;
	    RECT 15.6000 13.6000 16.4000 14.4000 ;
	    RECT 9.3000 10.4000 9.9000 13.6000 ;
	    RECT 9.2000 9.6000 10.0000 10.4000 ;
         LAYER metal3 ;
	    RECT 9.2000 14.3000 10.0000 14.4000 ;
	    RECT 15.6000 14.3000 16.4000 14.4000 ;
	    RECT 9.2000 13.7000 24.3000 14.3000 ;
	    RECT 9.2000 13.6000 10.0000 13.7000 ;
	    RECT 15.6000 13.6000 16.4000 13.7000 ;
      END
   END sel
   OBS
         LAYER metal1 ;
	    RECT 0.4000 20.4000 20.4000 21.6000 ;
	    RECT 2.8000 15.8000 3.6000 20.4000 ;
	    RECT 4.4000 15.2000 5.2000 19.8000 ;
	    RECT 6.0000 15.8000 6.8000 20.4000 ;
	    RECT 8.6000 16.4000 9.4000 19.8000 ;
	    RECT 7.6000 15.8000 9.4000 16.4000 ;
	    RECT 10.8000 15.8000 11.6000 19.8000 ;
	    RECT 12.4000 16.0000 13.2000 19.8000 ;
	    RECT 14.0000 16.6000 14.8000 20.4000 ;
	    RECT 15.6000 16.0000 16.4000 19.8000 ;
	    RECT 12.4000 15.8000 16.4000 16.0000 ;
	    RECT 3.0000 14.6000 5.2000 15.2000 ;
	    RECT 3.0000 11.6000 3.6000 14.6000 ;
	    RECT 4.4000 11.6000 5.2000 13.2000 ;
	    RECT 7.6000 12.3000 8.4000 15.8000 ;
	    RECT 11.0000 14.4000 11.6000 15.8000 ;
	    RECT 12.6000 15.4000 16.2000 15.8000 ;
	    RECT 10.8000 13.6000 13.4000 14.4000 ;
	    RECT 7.6000 11.7000 11.5000 12.3000 ;
	    RECT 2.4000 10.8000 3.6000 11.6000 ;
	    RECT 3.0000 10.2000 3.6000 10.8000 ;
	    RECT 3.0000 9.6000 5.2000 10.2000 ;
	    RECT 2.8000 1.6000 3.6000 9.0000 ;
	    RECT 4.4000 2.2000 5.2000 9.6000 ;
	    RECT 6.0000 1.6000 6.8000 6.2000 ;
	    RECT 7.6000 2.2000 8.4000 11.7000 ;
	    RECT 10.9000 10.4000 11.5000 11.7000 ;
	    RECT 10.8000 10.2000 11.6000 10.4000 ;
	    RECT 12.8000 10.2000 13.4000 13.6000 ;
	    RECT 14.0000 12.3000 14.8000 13.2000 ;
	    RECT 17.2000 12.3000 18.0000 19.8000 ;
	    RECT 18.8000 17.8000 19.6000 20.4000 ;
	    RECT 14.0000 11.7000 18.0000 12.3000 ;
	    RECT 14.0000 11.6000 14.8000 11.7000 ;
	    RECT 10.8000 9.6000 12.2000 10.2000 ;
	    RECT 12.8000 9.6000 13.8000 10.2000 ;
	    RECT 11.6000 8.4000 12.2000 9.6000 ;
	    RECT 11.6000 7.6000 12.4000 8.4000 ;
	    RECT 9.2000 1.6000 10.0000 6.2000 ;
	    RECT 11.4000 1.6000 12.2000 6.2000 ;
	    RECT 13.0000 2.2000 13.8000 9.6000 ;
	    RECT 15.6000 1.6000 16.4000 10.2000 ;
	    RECT 17.2000 2.2000 18.0000 11.7000 ;
	    RECT 18.8000 1.6000 19.6000 6.2000 ;
	    RECT 0.4000 0.4000 20.4000 1.6000 ;
         LAYER metal2 ;
	    RECT 10.8000 13.6000 11.6000 14.4000 ;
	    RECT 10.9000 12.4000 11.5000 13.6000 ;
	    RECT 4.4000 11.6000 5.2000 12.4000 ;
	    RECT 10.8000 11.6000 11.6000 12.4000 ;
         LAYER metal3 ;
	    RECT 4.4000 12.3000 5.2000 12.4000 ;
	    RECT 10.8000 12.3000 11.6000 12.4000 ;
	    RECT 4.4000 11.7000 11.6000 12.3000 ;
	    RECT 4.4000 11.6000 5.2000 11.7000 ;
	    RECT 10.8000 11.6000 11.6000 11.7000 ;
   END
END mux_using_if
