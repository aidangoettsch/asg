magic
tech scmos
magscale 1 2
timestamp 1593098107
<< metal1 >>
rect 1882 1814 1894 1816
rect 1867 1806 1869 1814
rect 1877 1806 1879 1814
rect 1887 1806 1889 1814
rect 1897 1806 1899 1814
rect 1907 1806 1909 1814
rect 1882 1804 1894 1806
rect 621 1777 684 1783
rect 2509 1757 2556 1763
rect 45 1717 60 1723
rect 77 1717 115 1723
rect 510 1717 540 1723
rect 733 1717 770 1723
rect 1565 1717 1580 1723
rect 1988 1717 2035 1723
rect 2477 1697 2499 1703
rect 138 1636 140 1644
rect 2452 1636 2454 1644
rect 666 1614 678 1616
rect 651 1606 653 1614
rect 661 1606 663 1614
rect 671 1606 673 1614
rect 681 1606 683 1614
rect 691 1606 693 1614
rect 666 1604 678 1606
rect 842 1576 844 1584
rect 2276 1576 2278 1584
rect 2301 1517 2316 1523
rect 2333 1517 2355 1523
rect 509 1497 531 1503
rect 781 1497 819 1503
rect 1092 1497 1122 1503
rect 2260 1497 2275 1503
rect 2356 1497 2371 1503
rect 429 1477 467 1483
rect 461 1457 467 1477
rect 989 1477 1027 1483
rect 2397 1477 2419 1483
rect 2525 1477 2556 1483
rect 941 1457 963 1463
rect 1882 1414 1894 1416
rect 1867 1406 1869 1414
rect 1877 1406 1879 1414
rect 1887 1406 1889 1414
rect 1897 1406 1899 1414
rect 1907 1406 1909 1414
rect 1882 1404 1894 1406
rect 637 1377 700 1383
rect 2202 1376 2204 1384
rect 1101 1357 1123 1363
rect 1988 1357 2028 1363
rect 2036 1357 2067 1363
rect 558 1337 588 1343
rect 1085 1337 1100 1343
rect 125 1317 163 1323
rect 1149 1317 1202 1323
rect 1965 1277 1980 1283
rect 186 1236 188 1244
rect 666 1214 678 1216
rect 651 1206 653 1214
rect 661 1206 663 1214
rect 671 1206 673 1214
rect 681 1206 683 1214
rect 691 1206 693 1214
rect 666 1204 678 1206
rect 2010 1176 2012 1184
rect 840 1136 844 1144
rect 1501 1097 1516 1103
rect 1725 1103 1731 1123
rect 1725 1097 1763 1103
rect 1773 1097 1820 1103
rect 1837 1097 1916 1103
rect 2420 1097 2451 1103
rect 740 1077 787 1083
rect 1661 1077 1692 1083
rect 2365 1057 2412 1063
rect 1882 1014 1894 1016
rect 1867 1006 1869 1014
rect 1877 1006 1879 1014
rect 1887 1006 1889 1014
rect 1897 1006 1899 1014
rect 1907 1006 1909 1014
rect 1882 1004 1894 1006
rect 616 976 620 984
rect 1805 977 1820 983
rect 477 957 499 963
rect 269 937 323 943
rect 548 937 563 943
rect 653 937 716 943
rect 125 917 163 923
rect 1092 917 1107 923
rect 1181 917 1220 923
rect 1212 916 1220 917
rect 1268 917 1283 923
rect 708 897 755 903
rect 1949 877 1964 883
rect 2525 877 2556 883
rect 186 836 188 844
rect 1108 836 1110 844
rect 666 814 678 816
rect 651 806 653 814
rect 661 806 663 814
rect 671 806 673 814
rect 681 806 683 814
rect 691 806 693 814
rect 666 804 678 806
rect 1668 776 1670 784
rect 1562 736 1564 744
rect 1021 697 1036 703
rect 1572 697 1619 703
rect 1629 697 1644 703
rect 1693 703 1699 723
rect 1693 697 1731 703
rect 1949 697 1987 703
rect 2397 697 2435 703
rect 1485 677 1500 683
rect 1757 677 1772 683
rect 1837 677 1932 683
rect 2541 677 2556 683
rect 717 657 764 663
rect 1853 657 1900 663
rect 2260 657 2275 663
rect 1882 614 1894 616
rect 1867 606 1869 614
rect 1877 606 1879 614
rect 1887 606 1889 614
rect 1897 606 1899 614
rect 1907 606 1909 614
rect 1882 604 1894 606
rect 2404 576 2406 584
rect 797 557 819 563
rect 1901 557 1980 563
rect 2436 557 2451 563
rect 740 537 771 543
rect 1924 537 2019 543
rect 2253 537 2291 543
rect 2324 537 2339 543
rect 45 517 60 523
rect 221 517 259 523
rect 317 517 332 523
rect 2285 517 2323 523
rect 1901 477 1964 483
rect 282 436 284 444
rect 666 414 678 416
rect 651 406 653 414
rect 661 406 663 414
rect 671 406 673 414
rect 681 406 683 414
rect 691 406 693 414
rect 666 404 678 406
rect 740 377 755 383
rect 2250 376 2252 384
rect 2372 376 2374 384
rect 1997 337 2100 343
rect 2500 336 2502 344
rect 2084 317 2099 323
rect 45 297 60 303
rect 77 297 92 303
rect 125 283 131 303
rect 573 297 611 303
rect 669 297 716 303
rect 781 297 835 303
rect 2253 297 2307 303
rect 2317 297 2332 303
rect 2340 297 2371 303
rect 2509 297 2556 303
rect 125 277 156 283
rect 820 277 835 283
rect 2333 277 2348 283
rect 109 257 124 263
rect 932 257 963 263
rect 1636 257 1651 263
rect 1997 257 2044 263
rect 1882 214 1894 216
rect 1867 206 1869 214
rect 1877 206 1879 214
rect 1887 206 1889 214
rect 1897 206 1899 214
rect 1907 206 1909 214
rect 1882 204 1894 206
rect 733 157 796 163
rect 2429 157 2451 163
rect 1646 137 1676 143
rect 2365 137 2396 143
rect 1837 117 1939 123
rect 1812 96 1820 104
rect 1837 97 1843 117
rect 2509 77 2556 83
rect 2180 56 2182 64
rect 666 14 678 16
rect 651 6 653 14
rect 661 6 663 14
rect 671 6 673 14
rect 681 6 683 14
rect 691 6 693 14
rect 666 4 678 6
<< m2contact >>
rect 1859 1806 1867 1814
rect 1869 1806 1877 1814
rect 1879 1806 1887 1814
rect 1889 1806 1897 1814
rect 1899 1806 1907 1814
rect 1909 1806 1917 1814
rect 572 1776 580 1784
rect 684 1776 692 1784
rect 700 1776 708 1784
rect 1532 1776 1540 1784
rect 2060 1776 2068 1784
rect 60 1756 68 1764
rect 348 1756 356 1764
rect 924 1756 932 1764
rect 1340 1756 1348 1764
rect 1580 1756 1588 1764
rect 1788 1756 1796 1764
rect 2236 1756 2244 1764
rect 2556 1756 2564 1764
rect 316 1736 324 1744
rect 956 1736 964 1744
rect 1100 1736 1108 1744
rect 1308 1736 1316 1744
rect 1820 1736 1828 1744
rect 2204 1736 2212 1744
rect 2428 1736 2436 1744
rect 60 1716 68 1724
rect 156 1716 164 1724
rect 172 1716 180 1724
rect 316 1716 324 1724
rect 540 1716 548 1724
rect 588 1716 596 1724
rect 1052 1716 1060 1724
rect 1196 1716 1204 1724
rect 1420 1716 1428 1724
rect 1580 1716 1588 1724
rect 1916 1716 1924 1724
rect 1980 1716 1988 1724
rect 2124 1716 2132 1724
rect 2444 1716 2452 1724
rect 220 1696 228 1704
rect 1052 1696 1060 1704
rect 1212 1696 1220 1704
rect 1916 1696 1924 1704
rect 2108 1696 2116 1704
rect 12 1676 20 1684
rect 140 1636 148 1644
rect 220 1636 228 1644
rect 764 1636 772 1644
rect 1052 1636 1060 1644
rect 1148 1636 1156 1644
rect 1212 1636 1220 1644
rect 1500 1636 1508 1644
rect 1596 1636 1604 1644
rect 1628 1636 1636 1644
rect 1916 1636 1924 1644
rect 2108 1636 2116 1644
rect 2396 1636 2404 1644
rect 2444 1636 2452 1644
rect 643 1606 651 1614
rect 653 1606 661 1614
rect 663 1606 671 1614
rect 673 1606 681 1614
rect 683 1606 691 1614
rect 693 1606 701 1614
rect 28 1576 36 1584
rect 316 1576 324 1584
rect 364 1576 372 1584
rect 460 1576 468 1584
rect 620 1576 628 1584
rect 844 1576 852 1584
rect 1052 1576 1060 1584
rect 1468 1576 1476 1584
rect 1756 1576 1764 1584
rect 1804 1576 1812 1584
rect 1916 1576 1924 1584
rect 2204 1576 2212 1584
rect 2268 1576 2276 1584
rect 1372 1558 1380 1566
rect 1020 1536 1028 1544
rect 2476 1536 2484 1544
rect 316 1516 324 1524
rect 940 1516 948 1524
rect 1372 1512 1380 1520
rect 1756 1516 1764 1524
rect 2204 1516 2212 1524
rect 2316 1516 2324 1524
rect 284 1496 292 1504
rect 396 1496 404 1504
rect 412 1496 420 1504
rect 588 1496 596 1504
rect 748 1496 756 1504
rect 860 1496 868 1504
rect 876 1496 884 1504
rect 908 1496 916 1504
rect 1004 1496 1012 1504
rect 1084 1496 1092 1504
rect 1404 1496 1412 1504
rect 1548 1496 1556 1504
rect 1996 1496 2004 1504
rect 2108 1496 2116 1504
rect 2252 1496 2260 1504
rect 2348 1496 2356 1504
rect 2380 1496 2388 1504
rect 2444 1496 2452 1504
rect 2492 1496 2500 1504
rect 220 1476 228 1484
rect 188 1456 196 1464
rect 444 1456 452 1464
rect 492 1476 500 1484
rect 556 1476 564 1484
rect 732 1476 740 1484
rect 892 1476 900 1484
rect 972 1476 980 1484
rect 1308 1476 1316 1484
rect 1660 1476 1668 1484
rect 2108 1476 2116 1484
rect 2252 1476 2260 1484
rect 2556 1476 2564 1484
rect 540 1456 548 1464
rect 572 1456 580 1464
rect 700 1456 708 1464
rect 764 1456 772 1464
rect 1036 1456 1044 1464
rect 1276 1456 1284 1464
rect 1628 1456 1636 1464
rect 1820 1456 1828 1464
rect 2076 1456 2084 1464
rect 2316 1456 2324 1464
rect 2428 1456 2436 1464
rect 716 1436 724 1444
rect 2412 1436 2420 1444
rect 1859 1406 1867 1414
rect 1869 1406 1877 1414
rect 1879 1406 1887 1414
rect 1889 1406 1897 1414
rect 1899 1406 1907 1414
rect 1909 1406 1917 1414
rect 700 1376 708 1384
rect 732 1376 740 1384
rect 1196 1376 1204 1384
rect 1564 1376 1572 1384
rect 1612 1376 1620 1384
rect 2204 1376 2212 1384
rect 2236 1376 2244 1384
rect 108 1356 116 1364
rect 396 1356 404 1364
rect 892 1356 900 1364
rect 1356 1356 1364 1364
rect 1628 1356 1636 1364
rect 1804 1356 1812 1364
rect 1980 1356 1988 1364
rect 2028 1356 2036 1364
rect 2492 1356 2500 1364
rect 12 1336 20 1344
rect 60 1336 68 1344
rect 364 1336 372 1344
rect 588 1336 596 1344
rect 924 1336 932 1344
rect 1100 1336 1108 1344
rect 1164 1336 1172 1344
rect 1388 1336 1396 1344
rect 1596 1336 1604 1344
rect 1772 1336 1780 1344
rect 2172 1336 2180 1344
rect 2204 1336 2212 1344
rect 2284 1336 2292 1344
rect 2316 1336 2324 1344
rect 2348 1336 2356 1344
rect 44 1316 52 1324
rect 92 1316 100 1324
rect 204 1316 212 1324
rect 220 1316 228 1324
rect 284 1316 292 1324
rect 476 1316 484 1324
rect 604 1316 612 1324
rect 812 1316 820 1324
rect 1020 1316 1028 1324
rect 1068 1316 1076 1324
rect 1484 1316 1492 1324
rect 1532 1316 1540 1324
rect 1580 1316 1588 1324
rect 1676 1316 1684 1324
rect 2076 1316 2084 1324
rect 2108 1316 2116 1324
rect 2156 1316 2164 1324
rect 2220 1316 2228 1324
rect 2268 1316 2276 1324
rect 2332 1316 2340 1324
rect 2380 1316 2388 1324
rect 2444 1316 2452 1324
rect 300 1300 308 1308
rect 636 1296 644 1304
rect 988 1300 996 1308
rect 1116 1296 1124 1304
rect 1452 1300 1460 1308
rect 1676 1296 1684 1304
rect 2092 1296 2100 1304
rect 2300 1296 2308 1304
rect 2364 1296 2372 1304
rect 2428 1296 2436 1304
rect 1980 1276 1988 1284
rect 2124 1276 2132 1284
rect 2396 1276 2404 1284
rect 2460 1276 2468 1284
rect 2508 1276 2516 1284
rect 300 1254 308 1262
rect 988 1254 996 1262
rect 1452 1254 1460 1262
rect 2380 1256 2388 1264
rect 2444 1256 2452 1264
rect 188 1236 196 1244
rect 556 1236 564 1244
rect 732 1236 740 1244
rect 1676 1236 1684 1244
rect 2108 1236 2116 1244
rect 643 1206 651 1214
rect 653 1206 661 1214
rect 663 1206 671 1214
rect 673 1206 681 1214
rect 683 1206 691 1214
rect 693 1206 701 1214
rect 28 1176 36 1184
rect 316 1176 324 1184
rect 396 1176 404 1184
rect 1020 1176 1028 1184
rect 1068 1176 1076 1184
rect 1228 1176 1236 1184
rect 1260 1176 1268 1184
rect 1436 1176 1444 1184
rect 1564 1176 1572 1184
rect 1708 1176 1716 1184
rect 1964 1176 1972 1184
rect 2012 1176 2020 1184
rect 2076 1176 2084 1184
rect 844 1136 852 1144
rect 1276 1136 1284 1144
rect 1580 1136 1588 1144
rect 1612 1136 1620 1144
rect 1740 1136 1748 1144
rect 1948 1136 1956 1144
rect 316 1116 324 1124
rect 396 1116 404 1124
rect 1004 1116 1012 1124
rect 1308 1116 1316 1124
rect 1548 1116 1556 1124
rect 284 1096 292 1104
rect 492 1096 500 1104
rect 892 1096 900 1104
rect 924 1096 932 1104
rect 972 1096 980 1104
rect 1052 1096 1060 1104
rect 1100 1096 1108 1104
rect 1292 1096 1300 1104
rect 1516 1096 1524 1104
rect 1564 1096 1572 1104
rect 1852 1116 1860 1124
rect 1980 1116 1988 1124
rect 2076 1116 2084 1124
rect 1820 1096 1828 1104
rect 1916 1096 1924 1104
rect 1964 1096 1972 1104
rect 1996 1096 2004 1104
rect 2076 1096 2084 1104
rect 2412 1096 2420 1104
rect 220 1076 228 1084
rect 492 1076 500 1084
rect 732 1076 740 1084
rect 876 1076 884 1084
rect 908 1076 916 1084
rect 956 1076 964 1084
rect 988 1076 996 1084
rect 1116 1076 1124 1084
rect 1324 1076 1332 1084
rect 1644 1076 1652 1084
rect 1692 1076 1700 1084
rect 1788 1076 1796 1084
rect 1804 1076 1812 1084
rect 2172 1076 2180 1084
rect 2444 1076 2452 1084
rect 188 1056 196 1064
rect 524 1056 532 1064
rect 940 1056 948 1064
rect 1516 1056 1524 1064
rect 1628 1056 1636 1064
rect 2028 1056 2036 1064
rect 2204 1056 2212 1064
rect 2412 1056 2420 1064
rect 684 1036 692 1044
rect 1020 1036 1028 1044
rect 1068 1036 1076 1044
rect 1468 1036 1476 1044
rect 1532 1036 1540 1044
rect 2428 1036 2436 1044
rect 1859 1006 1867 1014
rect 1869 1006 1877 1014
rect 1879 1006 1887 1014
rect 1889 1006 1897 1014
rect 1899 1006 1907 1014
rect 1909 1006 1917 1014
rect 332 976 340 984
rect 460 976 468 984
rect 620 976 628 984
rect 1308 976 1316 984
rect 1820 976 1828 984
rect 1996 976 2004 984
rect 2460 976 2468 984
rect 108 956 116 964
rect 236 956 244 964
rect 252 956 260 964
rect 284 956 292 964
rect 348 956 356 964
rect 908 956 916 964
rect 1484 956 1492 964
rect 1740 956 1748 964
rect 1916 956 1924 964
rect 2092 956 2100 964
rect 2300 956 2308 964
rect 12 936 20 944
rect 60 936 68 944
rect 364 936 372 944
rect 396 936 404 944
rect 444 936 452 944
rect 540 936 548 944
rect 716 936 724 944
rect 940 936 948 944
rect 1084 936 1092 944
rect 1148 936 1156 944
rect 1196 936 1204 944
rect 1452 936 1460 944
rect 1646 936 1654 944
rect 1676 936 1684 944
rect 1692 932 1700 940
rect 1964 936 1972 944
rect 2108 936 2116 944
rect 2268 936 2276 944
rect 44 916 52 924
rect 92 916 100 924
rect 204 916 212 924
rect 220 916 228 924
rect 268 916 276 924
rect 300 916 308 924
rect 380 916 388 924
rect 428 916 436 924
rect 524 916 532 924
rect 1020 916 1028 924
rect 1084 916 1092 924
rect 1244 916 1252 924
rect 1260 916 1268 924
rect 1372 916 1380 924
rect 1772 916 1780 924
rect 1820 916 1828 924
rect 1948 916 1956 924
rect 2044 916 2052 924
rect 2172 916 2180 924
rect 2492 916 2500 924
rect 412 896 420 904
rect 492 896 500 904
rect 700 896 708 904
rect 1004 900 1012 908
rect 1132 896 1140 904
rect 1388 900 1396 908
rect 1836 896 1844 904
rect 1996 896 2004 904
rect 2060 896 2068 904
rect 2204 900 2212 908
rect 1804 876 1812 884
rect 1964 876 1972 884
rect 2028 876 2036 884
rect 2556 876 2564 884
rect 2204 854 2212 862
rect 188 836 196 844
rect 1004 836 1012 844
rect 1100 836 1108 844
rect 1388 836 1396 844
rect 1724 836 1732 844
rect 1772 836 1780 844
rect 2044 836 2052 844
rect 2076 836 2084 844
rect 2124 836 2132 844
rect 2460 836 2468 844
rect 643 806 651 814
rect 653 806 661 814
rect 663 806 671 814
rect 673 806 681 814
rect 683 806 691 814
rect 693 806 701 814
rect 28 776 36 784
rect 316 776 324 784
rect 716 776 724 784
rect 860 776 868 784
rect 1116 776 1124 784
rect 1660 776 1668 784
rect 2060 776 2068 784
rect 2156 776 2164 784
rect 2380 776 2388 784
rect 460 758 468 766
rect 2476 756 2484 764
rect 1564 736 1572 744
rect 2076 736 2084 744
rect 2140 736 2148 744
rect 2172 736 2180 744
rect 316 716 324 724
rect 460 712 468 720
rect 924 716 932 724
rect 1116 716 1124 724
rect 1532 716 1540 724
rect 316 696 324 704
rect 428 696 436 704
rect 812 696 820 704
rect 892 696 900 704
rect 972 696 980 704
rect 1036 696 1044 704
rect 1116 696 1124 704
rect 1148 696 1156 704
rect 1468 696 1476 704
rect 1564 696 1572 704
rect 1644 696 1652 704
rect 1660 696 1668 704
rect 1708 716 1716 724
rect 1772 716 1780 724
rect 2012 716 2020 724
rect 2108 716 2116 724
rect 2204 716 2212 724
rect 2412 716 2420 724
rect 1740 696 1748 704
rect 1820 696 1828 704
rect 2028 696 2036 704
rect 2092 696 2100 704
rect 2188 696 2196 704
rect 2252 696 2260 704
rect 2332 696 2340 704
rect 2444 696 2452 704
rect 2508 696 2516 704
rect 220 676 228 684
rect 524 676 532 684
rect 828 676 836 684
rect 876 676 884 684
rect 940 676 948 684
rect 1068 676 1076 684
rect 1212 676 1220 684
rect 1500 676 1508 684
rect 1516 676 1524 684
rect 1580 676 1588 684
rect 1644 676 1652 684
rect 1772 676 1780 684
rect 1804 676 1812 684
rect 1932 676 1940 684
rect 1964 676 1972 684
rect 1996 676 2004 684
rect 2348 676 2356 684
rect 2380 676 2388 684
rect 2460 676 2468 684
rect 2556 676 2564 684
rect 188 656 196 664
rect 364 656 372 664
rect 556 656 564 664
rect 764 656 772 664
rect 860 656 868 664
rect 924 656 932 664
rect 1244 656 1252 664
rect 1404 656 1412 664
rect 1500 656 1508 664
rect 1596 656 1604 664
rect 1788 656 1796 664
rect 1900 656 1908 664
rect 1932 656 1940 664
rect 2044 656 2052 664
rect 2124 656 2132 664
rect 2220 656 2228 664
rect 2252 656 2260 664
rect 2284 656 2292 664
rect 2300 656 2308 664
rect 2492 656 2500 664
rect 380 636 388 644
rect 988 636 996 644
rect 1436 636 1444 644
rect 2236 636 2244 644
rect 2316 636 2324 644
rect 1859 606 1867 614
rect 1869 606 1877 614
rect 1879 606 1887 614
rect 1889 606 1897 614
rect 1899 606 1907 614
rect 1909 606 1917 614
rect 780 576 788 584
rect 892 576 900 584
rect 1548 576 1556 584
rect 2060 576 2068 584
rect 2348 576 2356 584
rect 2396 576 2404 584
rect 204 556 212 564
rect 508 556 516 564
rect 1068 556 1076 564
rect 1388 556 1396 564
rect 1740 556 1748 564
rect 1980 556 1988 564
rect 2076 556 2084 564
rect 2300 556 2308 564
rect 2364 556 2372 564
rect 2428 556 2436 564
rect 2460 556 2468 564
rect 60 536 68 544
rect 188 536 196 544
rect 540 536 548 544
rect 732 536 740 544
rect 860 536 868 544
rect 1004 536 1012 544
rect 1036 536 1044 544
rect 1084 536 1092 544
rect 1212 536 1220 544
rect 1356 536 1364 544
rect 1708 536 1716 544
rect 1916 536 1924 544
rect 2028 536 2036 544
rect 2092 536 2100 544
rect 2140 536 2148 544
rect 2316 536 2324 544
rect 2380 536 2388 544
rect 2508 536 2516 544
rect 60 516 68 524
rect 300 516 308 524
rect 332 516 340 524
rect 428 516 436 524
rect 748 516 756 524
rect 844 516 852 524
rect 1020 516 1028 524
rect 1468 516 1476 524
rect 1628 516 1636 524
rect 2044 516 2052 524
rect 2124 516 2132 524
rect 2156 516 2164 524
rect 2220 516 2228 524
rect 2236 516 2244 524
rect 2268 516 2276 524
rect 2428 516 2436 524
rect 636 496 644 504
rect 812 496 820 504
rect 1260 496 1268 504
rect 1644 500 1652 508
rect 1996 496 2004 504
rect 2092 496 2100 504
rect 2204 496 2212 504
rect 2412 496 2420 504
rect 2476 496 2484 504
rect 12 476 20 484
rect 1964 476 1972 484
rect 2188 476 2196 484
rect 1468 454 1476 462
rect 1644 454 1652 462
rect 284 436 292 444
rect 348 436 356 444
rect 636 436 644 444
rect 1068 436 1076 444
rect 1548 436 1556 444
rect 2492 436 2500 444
rect 643 406 651 414
rect 653 406 661 414
rect 663 406 671 414
rect 673 406 681 414
rect 683 406 691 414
rect 693 406 701 414
rect 220 376 228 384
rect 508 376 516 384
rect 620 376 628 384
rect 732 376 740 384
rect 1612 376 1620 384
rect 1660 376 1668 384
rect 1708 376 1716 384
rect 2252 376 2260 384
rect 2364 376 2372 384
rect 2428 376 2436 384
rect 1212 358 1220 366
rect 1356 358 1364 366
rect 12 336 20 344
rect 2444 336 2452 344
rect 2492 336 2500 344
rect 508 316 516 324
rect 1212 312 1220 320
rect 1356 312 1364 320
rect 1708 316 1716 324
rect 2076 316 2084 324
rect 2220 316 2228 324
rect 2284 316 2292 324
rect 2396 316 2404 324
rect 2412 316 2420 324
rect 60 296 68 304
rect 92 296 100 304
rect 140 296 148 304
rect 300 296 308 304
rect 476 296 484 304
rect 652 296 660 304
rect 716 296 724 304
rect 876 296 884 304
rect 892 296 900 304
rect 908 296 916 304
rect 1148 296 1156 304
rect 1260 296 1268 304
rect 1324 296 1332 304
rect 1532 296 1540 304
rect 1708 296 1716 304
rect 2124 296 2132 304
rect 2188 296 2196 304
rect 2332 296 2340 304
rect 2428 296 2436 304
rect 2556 296 2564 304
rect 156 276 164 284
rect 412 276 420 284
rect 812 276 820 284
rect 1148 276 1156 284
rect 1420 276 1428 284
rect 1804 276 1812 284
rect 2108 276 2116 284
rect 2140 276 2148 284
rect 2204 276 2212 284
rect 2268 276 2276 284
rect 2348 276 2356 284
rect 60 256 68 264
rect 92 256 100 264
rect 124 256 132 264
rect 188 256 196 264
rect 380 256 388 264
rect 556 256 564 264
rect 764 256 772 264
rect 796 256 804 264
rect 924 256 932 264
rect 1116 256 1124 264
rect 1452 256 1460 264
rect 1628 256 1636 264
rect 1836 256 1844 264
rect 2044 256 2052 264
rect 2476 256 2484 264
rect 172 236 180 244
rect 2156 236 2164 244
rect 1859 206 1867 214
rect 1869 206 1877 214
rect 1879 206 1887 214
rect 1889 206 1897 214
rect 1899 206 1907 214
rect 1909 206 1917 214
rect 28 176 36 184
rect 1292 176 1300 184
rect 2140 176 2148 184
rect 2332 176 2340 184
rect 2412 176 2420 184
rect 188 156 196 164
rect 572 156 580 164
rect 796 156 804 164
rect 1132 156 1140 164
rect 1484 156 1492 164
rect 1980 156 1988 164
rect 2220 156 2228 164
rect 2460 156 2468 164
rect 220 136 228 144
rect 540 136 548 144
rect 1100 136 1108 144
rect 1452 136 1460 144
rect 1676 136 1684 144
rect 1772 136 1780 144
rect 1788 136 1796 144
rect 1964 136 1972 144
rect 2012 136 2020 144
rect 2092 136 2100 144
rect 2156 136 2164 144
rect 2396 136 2404 144
rect 300 116 308 124
rect 396 116 404 124
rect 476 116 484 124
rect 652 116 660 124
rect 860 116 868 124
rect 876 116 884 124
rect 924 116 932 124
rect 1004 116 1012 124
rect 1356 116 1364 124
rect 1724 116 1732 124
rect 1804 116 1812 124
rect 284 100 292 108
rect 444 96 452 104
rect 1036 100 1044 108
rect 1388 100 1396 108
rect 1804 96 1812 104
rect 1948 116 1956 124
rect 2028 116 2036 124
rect 2044 116 2052 124
rect 2108 116 2116 124
rect 2172 116 2180 124
rect 2252 116 2260 124
rect 2300 116 2308 124
rect 2380 116 2388 124
rect 2476 116 2484 124
rect 1916 96 1924 104
rect 1980 96 1988 104
rect 2140 96 2148 104
rect 2236 96 2244 104
rect 2316 96 2324 104
rect 2332 96 2340 104
rect 2204 76 2212 84
rect 2284 76 2292 84
rect 2556 76 2564 84
rect 1036 54 1044 62
rect 2172 56 2180 64
rect 284 36 292 44
rect 364 36 372 44
rect 444 36 452 44
rect 828 36 836 44
rect 908 36 916 44
rect 956 36 964 44
rect 1388 36 1396 44
rect 2076 36 2084 44
rect 2268 36 2276 44
rect 643 6 651 14
rect 653 6 661 14
rect 663 6 671 14
rect 673 6 681 14
rect 683 6 691 14
rect 693 6 701 14
<< metal2 >>
rect 381 1824 387 1863
rect 557 1857 579 1863
rect 605 1857 627 1863
rect 573 1784 579 1857
rect 61 1724 67 1756
rect 13 1684 19 1696
rect 61 1604 67 1716
rect 173 1684 179 1716
rect 221 1644 227 1696
rect 141 1604 147 1636
rect 317 1624 323 1716
rect 29 1584 35 1596
rect 221 1484 227 1596
rect 285 1504 291 1616
rect 317 1524 323 1576
rect 189 1404 195 1456
rect 29 1357 44 1363
rect 29 1184 35 1357
rect 45 1324 51 1356
rect 61 1304 67 1336
rect 221 1324 227 1416
rect 285 1324 291 1496
rect 349 1484 355 1756
rect 365 1584 371 1636
rect 461 1584 467 1736
rect 573 1717 588 1723
rect 397 1364 403 1476
rect 413 1424 419 1496
rect 445 1464 451 1496
rect 493 1424 499 1476
rect 541 1464 547 1716
rect 557 1484 563 1716
rect 573 1464 579 1717
rect 621 1584 627 1857
rect 685 1784 691 1796
rect 701 1784 707 1816
rect 733 1804 739 1863
rect 765 1824 771 1863
rect 666 1614 678 1616
rect 651 1606 653 1614
rect 661 1606 663 1614
rect 671 1606 673 1614
rect 681 1606 683 1614
rect 691 1606 693 1614
rect 666 1604 678 1606
rect 573 1384 579 1456
rect 589 1344 595 1496
rect 93 1004 99 1316
rect 189 1084 195 1236
rect 285 1104 291 1316
rect 301 1262 307 1300
rect 365 1224 371 1336
rect 605 1324 611 1496
rect 301 1083 307 1196
rect 317 1124 323 1176
rect 285 1077 307 1083
rect 189 984 195 1056
rect 237 964 243 996
rect 285 964 291 1077
rect 333 984 339 1216
rect 397 1124 403 1176
rect 493 1104 499 1316
rect 637 1304 643 1516
rect 765 1464 771 1636
rect 845 1584 851 1736
rect 861 1504 867 1536
rect 701 1384 707 1456
rect 717 1344 723 1436
rect 877 1424 883 1496
rect 893 1464 899 1476
rect 925 1364 931 1756
rect 1053 1644 1059 1696
rect 1069 1623 1075 1863
rect 1133 1824 1139 1863
rect 1533 1857 1555 1863
rect 2045 1857 2067 1863
rect 1101 1744 1107 1816
rect 1533 1784 1539 1857
rect 1882 1814 1894 1816
rect 1867 1806 1869 1814
rect 1877 1806 1879 1814
rect 1887 1806 1889 1814
rect 1897 1806 1899 1814
rect 1907 1806 1909 1814
rect 1882 1804 1894 1806
rect 2061 1784 2067 1857
rect 1213 1644 1219 1696
rect 1309 1644 1315 1736
rect 1053 1617 1075 1623
rect 1053 1584 1059 1617
rect 557 1204 563 1236
rect 666 1214 678 1216
rect 651 1206 653 1214
rect 661 1206 663 1214
rect 671 1206 673 1214
rect 681 1206 683 1214
rect 691 1206 693 1214
rect 666 1204 678 1206
rect 733 1084 739 1236
rect 845 1104 851 1136
rect 925 1104 931 1316
rect 1005 1304 1011 1496
rect 1085 1484 1091 1496
rect 1037 1464 1043 1476
rect 989 1262 995 1300
rect 1021 1184 1027 1316
rect 1069 1184 1075 1296
rect 1005 1124 1011 1176
rect 1037 1097 1052 1103
rect 957 1084 963 1096
rect 493 1024 499 1076
rect 29 957 44 963
rect 29 784 35 957
rect 45 924 51 956
rect 349 944 355 956
rect 365 944 371 996
rect 461 984 467 1016
rect 525 984 531 1056
rect 621 984 627 1076
rect 685 1004 691 1036
rect 877 1004 883 1076
rect 941 1064 947 1076
rect 973 1064 979 1096
rect 445 944 451 956
rect 61 904 67 936
rect 221 924 227 936
rect 93 904 99 916
rect 189 684 195 836
rect 317 724 323 776
rect 61 544 67 556
rect 189 544 195 656
rect 13 484 19 496
rect 13 324 19 336
rect 61 264 67 296
rect 157 284 163 456
rect 189 304 195 536
rect 205 524 211 556
rect 333 524 339 936
rect 541 904 547 936
rect 365 664 371 896
rect 413 884 419 896
rect 493 884 499 896
rect 413 744 419 876
rect 666 814 678 816
rect 651 806 653 814
rect 661 806 663 814
rect 671 806 673 814
rect 681 806 683 814
rect 691 806 693 814
rect 666 804 678 806
rect 717 784 723 936
rect 861 784 867 816
rect 461 720 467 758
rect 381 644 387 656
rect 381 524 387 636
rect 429 524 435 696
rect 525 644 531 676
rect 765 664 771 676
rect 557 624 563 656
rect 509 564 515 616
rect 205 383 211 516
rect 333 464 339 516
rect 205 377 220 383
rect 93 264 99 276
rect 61 184 67 256
rect 173 204 179 236
rect 205 203 211 296
rect 285 284 291 436
rect 429 424 435 516
rect 477 304 483 416
rect 509 404 515 556
rect 509 324 515 376
rect 189 197 211 203
rect 189 164 195 197
rect 221 144 227 196
rect 301 124 307 296
rect 381 264 387 296
rect 397 124 403 196
rect 477 124 483 296
rect 557 204 563 256
rect 541 144 547 176
rect 573 164 579 396
rect 621 384 627 536
rect 637 444 643 496
rect 666 414 678 416
rect 651 406 653 414
rect 661 406 663 414
rect 671 406 673 414
rect 681 406 683 414
rect 691 406 693 414
rect 666 404 678 406
rect 653 304 659 376
rect 717 324 723 456
rect 733 384 739 536
rect 717 304 723 316
rect 765 264 771 656
rect 781 584 787 636
rect 797 503 803 736
rect 829 664 835 676
rect 845 524 851 696
rect 909 683 915 956
rect 941 824 947 936
rect 1021 924 1027 1036
rect 1005 844 1011 900
rect 925 724 931 736
rect 1037 704 1043 1097
rect 1069 923 1075 1036
rect 1085 944 1091 1476
rect 1117 1304 1123 1516
rect 1117 1124 1123 1296
rect 1101 1064 1107 1096
rect 1117 1044 1123 1076
rect 1069 917 1084 923
rect 941 684 947 696
rect 893 677 915 683
rect 893 644 899 677
rect 893 624 899 636
rect 893 584 899 616
rect 797 497 812 503
rect 861 384 867 536
rect 893 304 899 316
rect 653 124 659 156
rect 765 124 771 256
rect 797 164 803 256
rect 813 184 819 276
rect 925 264 931 376
rect 797 144 803 156
rect 861 124 867 136
rect 925 124 931 256
rect 989 164 995 636
rect 1005 544 1011 556
rect 1085 544 1091 816
rect 1101 564 1107 836
rect 1117 824 1123 1036
rect 1133 904 1139 1116
rect 1149 1104 1155 1636
rect 1341 1624 1347 1756
rect 1581 1724 1587 1756
rect 1277 1464 1283 1616
rect 1373 1520 1379 1558
rect 1421 1504 1427 1716
rect 1469 1584 1475 1596
rect 1309 1484 1315 1496
rect 1197 1384 1203 1456
rect 1165 1184 1171 1336
rect 1229 1184 1235 1236
rect 1261 1184 1267 1416
rect 1277 1364 1283 1456
rect 1277 1244 1283 1356
rect 1485 1324 1491 1336
rect 1453 1262 1459 1300
rect 1437 1184 1443 1216
rect 1197 944 1203 1176
rect 1277 1084 1283 1136
rect 1309 1124 1315 1156
rect 1293 1104 1299 1116
rect 1501 1083 1507 1636
rect 1581 1604 1587 1716
rect 1597 1604 1603 1636
rect 1757 1524 1763 1576
rect 1549 1423 1555 1496
rect 1661 1424 1667 1476
rect 1789 1464 1795 1756
rect 1821 1643 1827 1736
rect 1917 1644 1923 1696
rect 1805 1637 1827 1643
rect 1805 1584 1811 1637
rect 1981 1584 1987 1716
rect 2109 1644 2115 1696
rect 2125 1623 2131 1716
rect 2205 1624 2211 1736
rect 2109 1617 2131 1623
rect 1805 1444 1811 1456
rect 1549 1417 1571 1423
rect 1565 1384 1571 1417
rect 1613 1384 1619 1416
rect 1565 1364 1571 1376
rect 1645 1363 1651 1376
rect 1805 1364 1811 1436
rect 1882 1414 1894 1416
rect 1867 1406 1869 1414
rect 1877 1406 1879 1414
rect 1887 1406 1889 1414
rect 1897 1406 1899 1414
rect 1907 1406 1909 1414
rect 1882 1404 1894 1406
rect 1636 1357 1651 1363
rect 1565 1344 1571 1356
rect 1517 1317 1532 1323
rect 1517 1104 1523 1317
rect 1565 1317 1580 1323
rect 1565 1184 1571 1317
rect 1549 1084 1555 1116
rect 1501 1077 1516 1083
rect 1309 1064 1315 1076
rect 1149 924 1155 936
rect 1245 924 1251 1056
rect 1309 984 1315 1056
rect 1325 1044 1331 1076
rect 1517 1064 1523 1076
rect 1565 1064 1571 1096
rect 1629 1064 1635 1156
rect 1645 1084 1651 1357
rect 1677 1324 1683 1356
rect 1677 1244 1683 1296
rect 1709 1184 1715 1336
rect 1805 1224 1811 1356
rect 1741 1144 1747 1176
rect 1949 1144 1955 1456
rect 1981 1364 1987 1576
rect 2109 1504 2115 1617
rect 2205 1524 2211 1576
rect 1965 1184 1971 1316
rect 1981 1184 1987 1276
rect 1997 1163 2003 1496
rect 2077 1444 2083 1456
rect 2013 1184 2019 1256
rect 1997 1157 2019 1163
rect 1693 1084 1699 1116
rect 1469 1004 1475 1036
rect 1533 1004 1539 1036
rect 1645 1003 1651 1076
rect 1629 997 1651 1003
rect 1373 924 1379 996
rect 1252 917 1260 923
rect 1117 724 1123 776
rect 1133 744 1139 896
rect 1117 684 1123 696
rect 1037 304 1043 536
rect 1069 404 1075 436
rect 1117 264 1123 636
rect 1149 304 1155 696
rect 1213 684 1219 736
rect 1245 704 1251 916
rect 1453 904 1459 936
rect 1389 844 1395 900
rect 1469 664 1475 696
rect 1245 644 1251 656
rect 1485 644 1491 956
rect 1501 684 1507 696
rect 1437 604 1443 636
rect 1213 544 1219 556
rect 1357 544 1363 596
rect 1213 320 1219 358
rect 1261 304 1267 496
rect 1389 404 1395 556
rect 1469 462 1475 516
rect 1357 320 1363 358
rect 1293 184 1299 276
rect 989 123 995 156
rect 989 117 1004 123
rect 285 44 291 100
rect 445 44 451 96
rect 1037 62 1043 100
rect 365 -17 371 36
rect 666 14 678 16
rect 651 6 653 14
rect 661 6 663 14
rect 671 6 673 14
rect 681 6 683 14
rect 691 6 693 14
rect 666 4 678 6
rect 829 -17 835 36
rect 909 -17 915 36
rect 957 -17 963 36
rect 365 -23 387 -17
rect 829 -23 851 -17
rect 893 -23 915 -17
rect 941 -23 963 -17
rect 1101 -17 1107 136
rect 1325 124 1331 296
rect 1453 264 1459 396
rect 1453 164 1459 256
rect 1549 204 1555 436
rect 1597 383 1603 656
rect 1629 584 1635 997
rect 1677 944 1683 1056
rect 1693 1003 1699 1076
rect 1805 1064 1811 1076
rect 1693 997 1715 1003
rect 1661 784 1667 896
rect 1661 704 1667 756
rect 1709 724 1715 997
rect 1741 944 1747 956
rect 1773 924 1779 1056
rect 1821 984 1827 1096
rect 1853 1084 1859 1116
rect 1882 1014 1894 1016
rect 1867 1006 1869 1014
rect 1877 1006 1879 1014
rect 1887 1006 1889 1014
rect 1897 1006 1899 1014
rect 1907 1006 1909 1014
rect 1882 1004 1894 1006
rect 1821 904 1827 916
rect 1837 904 1843 916
rect 1709 684 1715 716
rect 1725 703 1731 836
rect 1773 724 1779 836
rect 1773 704 1779 716
rect 1725 697 1740 703
rect 1773 684 1779 696
rect 1837 644 1843 896
rect 1901 684 1907 696
rect 1917 684 1923 956
rect 1949 924 1955 936
rect 1965 924 1971 936
rect 1965 884 1971 896
rect 1981 724 1987 1116
rect 1997 984 2003 1096
rect 2013 1044 2019 1157
rect 2029 1084 2035 1356
rect 2045 944 2051 1416
rect 2109 1404 2115 1476
rect 2084 1317 2108 1323
rect 2157 1304 2163 1316
rect 2093 1184 2099 1296
rect 2125 1264 2131 1276
rect 2173 1264 2179 1336
rect 2061 904 2067 1176
rect 2077 1124 2083 1176
rect 2109 1144 2115 1236
rect 2189 1183 2195 1436
rect 2205 1384 2211 1496
rect 2237 1444 2243 1756
rect 2269 1584 2275 1616
rect 2317 1504 2323 1516
rect 2237 1384 2243 1396
rect 2253 1384 2259 1476
rect 2285 1324 2291 1336
rect 2221 1284 2227 1316
rect 2269 1264 2275 1316
rect 2301 1304 2307 1376
rect 2317 1344 2323 1456
rect 2333 1324 2339 1716
rect 2429 1704 2435 1736
rect 2349 1344 2355 1356
rect 2365 1323 2371 1516
rect 2397 1484 2403 1636
rect 2429 1464 2435 1696
rect 2445 1524 2451 1636
rect 2557 1604 2563 1756
rect 2445 1484 2451 1496
rect 2365 1317 2380 1323
rect 2333 1204 2339 1316
rect 2413 1303 2419 1436
rect 2429 1364 2435 1456
rect 2413 1297 2428 1303
rect 2461 1284 2467 1496
rect 2493 1424 2499 1496
rect 2557 1484 2563 1496
rect 2397 1264 2403 1276
rect 2189 1177 2211 1183
rect 2077 1044 2083 1096
rect 2093 964 2099 1096
rect 2205 1064 2211 1177
rect 2413 1104 2419 1276
rect 2493 1204 2499 1356
rect 2029 884 2035 896
rect 1940 677 1964 683
rect 1901 664 1907 676
rect 1882 614 1894 616
rect 1867 606 1869 614
rect 1877 606 1879 614
rect 1887 606 1889 614
rect 1897 606 1899 614
rect 1907 606 1909 614
rect 1882 604 1894 606
rect 1597 377 1612 383
rect 1629 304 1635 516
rect 1645 462 1651 500
rect 1661 384 1667 416
rect 1709 324 1715 376
rect 1629 264 1635 276
rect 1677 144 1683 236
rect 1773 144 1779 156
rect 1789 144 1795 196
rect 1805 184 1811 276
rect 1837 264 1843 556
rect 1933 304 1939 656
rect 1981 564 1987 676
rect 1997 504 2003 676
rect 2013 504 2019 716
rect 2045 703 2051 836
rect 2061 784 2067 856
rect 2077 744 2083 836
rect 2045 697 2067 703
rect 2045 664 2051 676
rect 2061 664 2067 697
rect 2125 683 2131 836
rect 2157 784 2163 1016
rect 2173 924 2179 1036
rect 2205 964 2211 1056
rect 2205 862 2211 900
rect 2253 704 2259 736
rect 2109 677 2131 683
rect 2061 584 2067 636
rect 1882 214 1894 216
rect 1867 206 1869 214
rect 1877 206 1879 214
rect 1887 206 1889 214
rect 1897 206 1899 214
rect 1907 206 1909 214
rect 1882 204 1894 206
rect 1933 164 1939 296
rect 1965 224 1971 476
rect 1981 164 1987 496
rect 2077 324 2083 556
rect 2109 523 2115 677
rect 2189 664 2195 696
rect 2125 544 2131 656
rect 2269 643 2275 936
rect 2381 784 2387 1076
rect 2413 924 2419 1056
rect 2413 724 2419 916
rect 2429 884 2435 1036
rect 2445 1003 2451 1076
rect 2445 997 2467 1003
rect 2461 984 2467 997
rect 2557 884 2563 896
rect 2285 664 2291 696
rect 2253 637 2275 643
rect 2141 544 2147 556
rect 2109 517 2124 523
rect 1965 144 1971 156
rect 2013 144 2019 156
rect 1453 104 1459 136
rect 2013 104 2019 136
rect 2045 124 2051 256
rect 2093 144 2099 496
rect 2125 324 2131 516
rect 2141 284 2147 516
rect 2173 343 2179 536
rect 2237 524 2243 636
rect 2173 337 2195 343
rect 2141 244 2147 276
rect 2157 164 2163 236
rect 2109 124 2115 156
rect 2157 104 2163 136
rect 2173 124 2179 316
rect 2189 304 2195 337
rect 2221 324 2227 516
rect 2253 384 2259 637
rect 2269 544 2275 616
rect 2285 563 2291 656
rect 2317 644 2323 716
rect 2285 557 2300 563
rect 2317 544 2323 636
rect 2333 544 2339 696
rect 2356 677 2371 683
rect 2349 584 2355 636
rect 2365 584 2371 677
rect 2381 644 2387 676
rect 2413 664 2419 716
rect 2461 704 2467 836
rect 2445 624 2451 696
rect 2461 684 2467 696
rect 2557 684 2563 696
rect 2493 604 2499 656
rect 2461 564 2467 596
rect 2365 544 2371 556
rect 2509 544 2515 596
rect 2269 524 2275 536
rect 2285 324 2291 536
rect 2365 384 2371 496
rect 2381 464 2387 536
rect 2429 524 2435 536
rect 2477 504 2483 536
rect 2429 384 2435 456
rect 2493 364 2499 436
rect 2413 324 2419 356
rect 2269 204 2275 276
rect 2221 104 2227 156
rect 2285 144 2291 316
rect 2397 304 2403 316
rect 2333 184 2339 296
rect 2349 264 2355 276
rect 2413 223 2419 316
rect 2397 217 2419 223
rect 2301 124 2307 176
rect 2397 144 2403 217
rect 2413 184 2419 196
rect 1389 44 1395 100
rect 1101 -23 1139 -17
rect 2013 -23 2019 96
rect 2141 44 2147 96
rect 2253 84 2259 116
rect 2317 104 2323 136
rect 2381 104 2387 116
rect 2429 104 2435 296
rect 2461 164 2467 256
rect 2477 124 2483 216
rect 2557 84 2563 96
rect 2077 -17 2083 36
rect 2061 -23 2083 -17
rect 2205 -23 2211 76
rect 2285 64 2291 76
<< m3contact >>
rect 380 1816 388 1824
rect 316 1736 324 1744
rect 156 1716 164 1724
rect 12 1696 20 1704
rect 172 1676 180 1684
rect 284 1616 292 1624
rect 316 1616 324 1624
rect 28 1596 36 1604
rect 60 1596 68 1604
rect 140 1596 148 1604
rect 220 1596 228 1604
rect 220 1416 228 1424
rect 188 1396 196 1404
rect 12 1336 20 1344
rect 44 1356 52 1364
rect 108 1356 116 1364
rect 460 1736 468 1744
rect 364 1636 372 1644
rect 556 1716 564 1724
rect 396 1496 404 1504
rect 444 1496 452 1504
rect 348 1476 356 1484
rect 396 1476 404 1484
rect 444 1456 452 1464
rect 556 1476 564 1484
rect 700 1816 708 1824
rect 684 1796 692 1804
rect 764 1816 772 1824
rect 732 1796 740 1804
rect 844 1736 852 1744
rect 643 1606 651 1614
rect 653 1606 661 1614
rect 663 1606 671 1614
rect 673 1606 681 1614
rect 683 1606 691 1614
rect 693 1606 701 1614
rect 636 1516 644 1524
rect 604 1496 612 1504
rect 412 1416 420 1424
rect 492 1416 500 1424
rect 572 1376 580 1384
rect 396 1356 404 1364
rect 204 1316 212 1324
rect 60 1296 68 1304
rect 476 1316 484 1324
rect 492 1316 500 1324
rect 332 1216 340 1224
rect 364 1216 372 1224
rect 300 1196 308 1204
rect 188 1076 196 1084
rect 220 1076 228 1084
rect 92 996 100 1004
rect 236 996 244 1004
rect 188 976 196 984
rect 748 1496 756 1504
rect 732 1476 740 1484
rect 860 1536 868 1544
rect 908 1496 916 1504
rect 892 1456 900 1464
rect 876 1416 884 1424
rect 732 1376 740 1384
rect 956 1736 964 1744
rect 1052 1716 1060 1724
rect 1100 1816 1108 1824
rect 1132 1816 1140 1824
rect 1859 1806 1867 1814
rect 1869 1806 1877 1814
rect 1879 1806 1887 1814
rect 1889 1806 1897 1814
rect 1899 1806 1907 1814
rect 1909 1806 1917 1814
rect 1196 1716 1204 1724
rect 1308 1636 1316 1644
rect 1020 1536 1028 1544
rect 940 1516 948 1524
rect 1116 1516 1124 1524
rect 1004 1496 1012 1504
rect 972 1476 980 1484
rect 892 1356 900 1364
rect 924 1356 932 1364
rect 716 1336 724 1344
rect 924 1336 932 1344
rect 812 1316 820 1324
rect 924 1316 932 1324
rect 643 1206 651 1214
rect 653 1206 661 1214
rect 663 1206 671 1214
rect 673 1206 681 1214
rect 683 1206 691 1214
rect 693 1206 701 1214
rect 556 1196 564 1204
rect 1036 1476 1044 1484
rect 1084 1476 1092 1484
rect 1068 1316 1076 1324
rect 1004 1296 1012 1304
rect 1068 1296 1076 1304
rect 1004 1176 1012 1184
rect 844 1096 852 1104
rect 892 1096 900 1104
rect 956 1096 964 1104
rect 620 1076 628 1084
rect 908 1076 916 1084
rect 940 1076 948 1084
rect 460 1016 468 1024
rect 492 1016 500 1024
rect 364 996 372 1004
rect 12 936 20 944
rect 44 956 52 964
rect 108 956 116 964
rect 252 956 260 964
rect 988 1076 996 1084
rect 972 1056 980 1064
rect 684 996 692 1004
rect 876 996 884 1004
rect 524 976 532 984
rect 444 956 452 964
rect 220 936 228 944
rect 332 936 340 944
rect 348 936 356 944
rect 396 936 404 944
rect 204 916 212 924
rect 268 916 276 924
rect 300 916 308 924
rect 60 896 68 904
rect 92 896 100 904
rect 316 696 324 704
rect 188 676 196 684
rect 220 676 228 684
rect 188 656 196 664
rect 60 556 68 564
rect 60 516 68 524
rect 12 496 20 504
rect 156 456 164 464
rect 12 316 20 324
rect 92 296 100 304
rect 140 296 148 304
rect 380 916 388 924
rect 428 916 436 924
rect 524 916 532 924
rect 364 896 372 904
rect 540 896 548 904
rect 700 896 708 904
rect 412 876 420 884
rect 492 876 500 884
rect 643 806 651 814
rect 653 806 661 814
rect 663 806 671 814
rect 673 806 681 814
rect 683 806 691 814
rect 693 806 701 814
rect 860 816 868 824
rect 412 736 420 744
rect 796 736 804 744
rect 428 696 436 704
rect 380 656 388 664
rect 764 676 772 684
rect 524 636 532 644
rect 508 616 516 624
rect 556 616 564 624
rect 204 516 212 524
rect 300 516 308 524
rect 380 516 388 524
rect 332 456 340 464
rect 348 436 356 444
rect 188 296 196 304
rect 204 296 212 304
rect 92 276 100 284
rect 124 256 132 264
rect 188 256 196 264
rect 172 196 180 204
rect 428 416 436 424
rect 476 416 484 424
rect 540 536 548 544
rect 620 536 628 544
rect 508 396 516 404
rect 572 396 580 404
rect 380 296 388 304
rect 284 276 292 284
rect 28 176 36 184
rect 60 176 68 184
rect 220 196 228 204
rect 412 276 420 284
rect 396 196 404 204
rect 556 196 564 204
rect 540 176 548 184
rect 716 456 724 464
rect 643 406 651 414
rect 653 406 661 414
rect 663 406 671 414
rect 673 406 681 414
rect 683 406 691 414
rect 693 406 701 414
rect 652 376 660 384
rect 748 516 756 524
rect 732 376 740 384
rect 716 316 724 324
rect 780 636 788 644
rect 812 696 820 704
rect 844 696 852 704
rect 892 696 900 704
rect 828 656 836 664
rect 876 676 884 684
rect 940 816 948 824
rect 924 736 932 744
rect 1052 1096 1060 1104
rect 1100 1336 1108 1344
rect 1116 1116 1124 1124
rect 1132 1116 1140 1124
rect 1100 1056 1108 1064
rect 1116 1036 1124 1044
rect 1084 816 1092 824
rect 940 696 948 704
rect 972 696 980 704
rect 860 656 868 664
rect 1068 676 1076 684
rect 924 656 932 664
rect 892 636 900 644
rect 892 616 900 624
rect 844 516 852 524
rect 860 376 868 384
rect 924 376 932 384
rect 892 316 900 324
rect 876 296 884 304
rect 908 296 916 304
rect 652 156 660 164
rect 812 176 820 184
rect 796 136 804 144
rect 860 136 868 144
rect 1004 556 1012 564
rect 1068 556 1076 564
rect 1276 1616 1284 1624
rect 1340 1616 1348 1624
rect 1468 1596 1476 1604
rect 1308 1496 1316 1504
rect 1404 1496 1412 1504
rect 1420 1496 1428 1504
rect 1196 1456 1204 1464
rect 1260 1416 1268 1424
rect 1228 1236 1236 1244
rect 1276 1356 1284 1364
rect 1356 1356 1364 1364
rect 1388 1336 1396 1344
rect 1484 1336 1492 1344
rect 1276 1236 1284 1244
rect 1436 1216 1444 1224
rect 1164 1176 1172 1184
rect 1196 1176 1204 1184
rect 1148 1096 1156 1104
rect 1308 1156 1316 1164
rect 1292 1116 1300 1124
rect 1276 1076 1284 1084
rect 1308 1076 1316 1084
rect 1628 1636 1636 1644
rect 1580 1596 1588 1604
rect 1596 1596 1604 1604
rect 1548 1496 1556 1504
rect 1628 1456 1636 1464
rect 1916 1716 1924 1724
rect 2124 1716 2132 1724
rect 1916 1576 1924 1584
rect 1980 1576 1988 1584
rect 1788 1456 1796 1464
rect 1804 1456 1812 1464
rect 1820 1456 1828 1464
rect 1948 1456 1956 1464
rect 1804 1436 1812 1444
rect 1612 1416 1620 1424
rect 1660 1416 1668 1424
rect 1644 1376 1652 1384
rect 1564 1356 1572 1364
rect 1859 1406 1867 1414
rect 1869 1406 1877 1414
rect 1879 1406 1887 1414
rect 1889 1406 1897 1414
rect 1899 1406 1907 1414
rect 1909 1406 1917 1414
rect 1564 1336 1572 1344
rect 1596 1336 1604 1344
rect 1628 1156 1636 1164
rect 1580 1136 1588 1144
rect 1612 1136 1620 1144
rect 1516 1096 1524 1104
rect 1516 1076 1524 1084
rect 1548 1076 1556 1084
rect 1244 1056 1252 1064
rect 1308 1056 1316 1064
rect 1676 1356 1684 1364
rect 1708 1336 1716 1344
rect 1772 1336 1780 1344
rect 1804 1216 1812 1224
rect 1740 1176 1748 1184
rect 2204 1616 2212 1624
rect 2204 1496 2212 1504
rect 1964 1316 1972 1324
rect 1980 1176 1988 1184
rect 2076 1436 2084 1444
rect 2044 1416 2052 1424
rect 2012 1256 2020 1264
rect 1948 1136 1956 1144
rect 1692 1116 1700 1124
rect 1788 1076 1796 1084
rect 1564 1056 1572 1064
rect 1324 1036 1332 1044
rect 1468 1036 1476 1044
rect 1372 996 1380 1004
rect 1468 996 1476 1004
rect 1532 996 1540 1004
rect 1676 1056 1684 1064
rect 1148 916 1156 924
rect 1116 816 1124 824
rect 1132 736 1140 744
rect 1212 736 1220 744
rect 1116 676 1124 684
rect 1116 636 1124 644
rect 1100 556 1108 564
rect 1004 536 1012 544
rect 1084 536 1092 544
rect 1020 516 1028 524
rect 1068 396 1076 404
rect 1036 296 1044 304
rect 1452 896 1460 904
rect 1244 696 1252 704
rect 1404 656 1412 664
rect 1468 656 1476 664
rect 1564 736 1572 744
rect 1532 716 1540 724
rect 1500 696 1508 704
rect 1564 696 1572 704
rect 1516 676 1524 684
rect 1580 676 1588 684
rect 1500 656 1508 664
rect 1244 636 1252 644
rect 1484 636 1492 644
rect 1356 596 1364 604
rect 1436 596 1444 604
rect 1212 556 1220 564
rect 1548 576 1556 584
rect 1388 556 1396 564
rect 1388 396 1396 404
rect 1452 396 1460 404
rect 1260 296 1268 304
rect 1324 296 1332 304
rect 1148 276 1156 284
rect 1292 276 1300 284
rect 988 156 996 164
rect 1132 156 1140 164
rect 764 116 772 124
rect 876 116 884 124
rect 643 6 651 14
rect 653 6 661 14
rect 663 6 671 14
rect 673 6 681 14
rect 683 6 691 14
rect 693 6 701 14
rect 1420 276 1428 284
rect 1532 296 1540 304
rect 1772 1056 1780 1064
rect 1804 1056 1812 1064
rect 1644 936 1646 944
rect 1646 936 1652 944
rect 1692 940 1700 944
rect 1692 936 1700 940
rect 1660 896 1668 904
rect 1660 756 1668 764
rect 1740 936 1748 944
rect 1916 1096 1924 1104
rect 1964 1096 1972 1104
rect 1852 1076 1860 1084
rect 1859 1006 1867 1014
rect 1869 1006 1877 1014
rect 1879 1006 1887 1014
rect 1889 1006 1897 1014
rect 1899 1006 1907 1014
rect 1909 1006 1917 1014
rect 1836 916 1844 924
rect 1820 896 1828 904
rect 1804 876 1812 884
rect 1708 716 1716 724
rect 1644 696 1652 704
rect 1772 696 1780 704
rect 1820 696 1828 704
rect 1644 676 1652 684
rect 1708 676 1716 684
rect 1804 676 1812 684
rect 1788 656 1796 664
rect 1900 696 1908 704
rect 1948 936 1956 944
rect 1964 916 1972 924
rect 1964 896 1972 904
rect 2028 1076 2036 1084
rect 2028 1056 2036 1064
rect 2012 1036 2020 1044
rect 2188 1436 2196 1444
rect 2108 1396 2116 1404
rect 2092 1296 2100 1304
rect 2156 1296 2164 1304
rect 2124 1256 2132 1264
rect 2172 1256 2180 1264
rect 2060 1176 2068 1184
rect 2092 1176 2100 1184
rect 2044 936 2052 944
rect 2044 916 2052 924
rect 2332 1716 2340 1724
rect 2268 1616 2276 1624
rect 2252 1496 2260 1504
rect 2316 1496 2324 1504
rect 2236 1436 2244 1444
rect 2236 1396 2244 1404
rect 2252 1376 2260 1384
rect 2300 1376 2308 1384
rect 2204 1336 2212 1344
rect 2284 1316 2292 1324
rect 2220 1276 2228 1284
rect 2444 1716 2452 1724
rect 2428 1696 2436 1704
rect 2364 1516 2372 1524
rect 2348 1496 2356 1504
rect 2348 1356 2356 1364
rect 2380 1496 2388 1504
rect 2396 1476 2404 1484
rect 2556 1596 2564 1604
rect 2476 1536 2484 1544
rect 2444 1516 2452 1524
rect 2460 1496 2468 1504
rect 2556 1496 2564 1504
rect 2444 1476 2452 1484
rect 2300 1296 2308 1304
rect 2268 1256 2276 1264
rect 2364 1296 2372 1304
rect 2428 1356 2436 1364
rect 2444 1316 2452 1324
rect 2492 1416 2500 1424
rect 2412 1276 2420 1284
rect 2460 1276 2468 1284
rect 2380 1256 2388 1264
rect 2396 1256 2404 1264
rect 2332 1196 2340 1204
rect 2108 1136 2116 1144
rect 2092 1096 2100 1104
rect 2076 1036 2084 1044
rect 2172 1076 2180 1084
rect 2444 1256 2452 1264
rect 2508 1276 2516 1284
rect 2492 1196 2500 1204
rect 2412 1096 2420 1104
rect 2380 1076 2388 1084
rect 2172 1036 2180 1044
rect 2156 1016 2164 1024
rect 2108 936 2116 944
rect 1996 896 2004 904
rect 2028 896 2036 904
rect 2060 856 2068 864
rect 1980 716 1988 724
rect 2012 716 2020 724
rect 1900 676 1908 684
rect 1916 676 1924 684
rect 1980 676 1988 684
rect 1932 656 1940 664
rect 1836 636 1844 644
rect 1859 606 1867 614
rect 1869 606 1877 614
rect 1879 606 1887 614
rect 1889 606 1897 614
rect 1899 606 1907 614
rect 1909 606 1917 614
rect 1628 576 1636 584
rect 1740 556 1748 564
rect 1836 556 1844 564
rect 1708 536 1716 544
rect 1660 416 1668 424
rect 1628 296 1636 304
rect 1708 296 1716 304
rect 1628 276 1636 284
rect 1676 236 1684 244
rect 1548 196 1556 204
rect 1452 156 1460 164
rect 1484 156 1492 164
rect 1788 196 1796 204
rect 1772 156 1780 164
rect 1916 536 1924 544
rect 2028 696 2036 704
rect 2108 716 2116 724
rect 2044 676 2052 684
rect 2092 696 2100 704
rect 2204 956 2212 964
rect 2300 956 2308 964
rect 2140 736 2148 744
rect 2172 736 2180 744
rect 2252 736 2260 744
rect 2204 716 2212 724
rect 2188 696 2196 704
rect 2060 656 2068 664
rect 2060 636 2068 644
rect 2028 536 2036 544
rect 2044 516 2052 524
rect 1980 496 1988 504
rect 2012 496 2020 504
rect 1932 296 1940 304
rect 1859 206 1867 214
rect 1869 206 1877 214
rect 1879 206 1887 214
rect 1889 206 1897 214
rect 1899 206 1907 214
rect 1909 206 1917 214
rect 1804 176 1812 184
rect 1964 216 1972 224
rect 2092 536 2100 544
rect 2124 656 2132 664
rect 2188 656 2196 664
rect 2220 656 2228 664
rect 2252 656 2260 664
rect 2412 916 2420 924
rect 2492 916 2500 924
rect 2556 896 2564 904
rect 2428 876 2436 884
rect 2316 716 2324 724
rect 2284 696 2292 704
rect 2300 656 2308 664
rect 2140 556 2148 564
rect 2124 536 2132 544
rect 2172 536 2180 544
rect 2140 516 2148 524
rect 2156 516 2164 524
rect 1932 156 1940 164
rect 1964 156 1972 164
rect 2012 156 2020 164
rect 1788 136 1796 144
rect 1324 116 1332 124
rect 1356 116 1364 124
rect 1724 116 1732 124
rect 1804 116 1812 124
rect 1948 116 1956 124
rect 2124 316 2132 324
rect 2124 296 2132 304
rect 2204 496 2212 504
rect 2188 476 2196 484
rect 2172 316 2180 324
rect 2108 276 2116 284
rect 2140 236 2148 244
rect 2140 176 2148 184
rect 2108 156 2116 164
rect 2156 156 2164 164
rect 2092 136 2100 144
rect 2028 116 2036 124
rect 2268 616 2276 624
rect 2348 636 2356 644
rect 2476 756 2484 764
rect 2460 696 2468 704
rect 2508 696 2516 704
rect 2556 696 2564 704
rect 2412 656 2420 664
rect 2380 636 2388 644
rect 2444 616 2452 624
rect 2460 596 2468 604
rect 2492 596 2500 604
rect 2508 596 2516 604
rect 2364 576 2372 584
rect 2396 576 2404 584
rect 2428 556 2436 564
rect 2268 536 2276 544
rect 2284 536 2292 544
rect 2332 536 2340 544
rect 2364 536 2372 544
rect 2428 536 2436 544
rect 2476 536 2484 544
rect 2364 496 2372 504
rect 2412 496 2420 504
rect 2380 456 2388 464
rect 2428 456 2436 464
rect 2412 356 2420 364
rect 2492 356 2500 364
rect 2444 336 2452 344
rect 2492 336 2500 344
rect 2204 276 2212 284
rect 2268 196 2276 204
rect 2172 116 2180 124
rect 2396 296 2404 304
rect 2348 256 2356 264
rect 2556 296 2564 304
rect 2300 176 2308 184
rect 2332 176 2340 184
rect 2284 136 2292 144
rect 2412 196 2420 204
rect 2316 136 2324 144
rect 1452 96 1460 104
rect 1804 96 1812 104
rect 1916 96 1924 104
rect 1980 96 1988 104
rect 2012 96 2020 104
rect 2156 96 2164 104
rect 2220 96 2228 104
rect 2236 96 2244 104
rect 2460 256 2468 264
rect 2476 256 2484 264
rect 2476 216 2484 224
rect 2332 96 2340 104
rect 2380 96 2388 104
rect 2428 96 2436 104
rect 2556 96 2564 104
rect 2204 76 2212 84
rect 2252 76 2260 84
rect 2172 56 2180 64
rect 2140 36 2148 44
rect 2284 56 2292 64
rect 2268 36 2276 44
<< metal3 >>
rect 372 1817 380 1823
rect 708 1817 764 1823
rect 1108 1817 1132 1823
rect 1858 1814 1918 1816
rect 1858 1806 1859 1814
rect 1868 1806 1869 1814
rect 1907 1806 1908 1814
rect 1917 1806 1918 1814
rect 1858 1804 1918 1806
rect 692 1797 732 1803
rect 324 1737 460 1743
rect 852 1737 956 1743
rect 164 1717 556 1723
rect 1060 1717 1196 1723
rect 1924 1717 2124 1723
rect 2340 1717 2444 1723
rect -35 1697 12 1703
rect 2436 1697 2595 1703
rect 180 1677 204 1683
rect 1316 1637 1580 1643
rect 1588 1637 1628 1643
rect 292 1617 316 1623
rect 1284 1617 1340 1623
rect 2212 1617 2268 1623
rect 642 1614 702 1616
rect 642 1606 643 1614
rect 652 1606 653 1614
rect 691 1606 692 1614
rect 701 1606 702 1614
rect 642 1604 702 1606
rect 36 1597 60 1603
rect 148 1597 220 1603
rect 1476 1597 1580 1603
rect 1604 1597 1612 1603
rect 2516 1597 2556 1603
rect 2564 1597 2595 1603
rect 1924 1577 1980 1583
rect 868 1537 1020 1543
rect 2484 1537 2595 1543
rect 644 1517 940 1523
rect 948 1517 1116 1523
rect 2372 1517 2444 1523
rect 404 1497 444 1503
rect 612 1497 748 1503
rect 756 1497 908 1503
rect 916 1497 1004 1503
rect 1021 1497 1308 1503
rect 356 1477 396 1483
rect 564 1477 732 1483
rect 1021 1483 1027 1497
rect 1412 1497 1420 1503
rect 1428 1497 1548 1503
rect 2212 1497 2252 1503
rect 2324 1497 2348 1503
rect 2388 1497 2460 1503
rect 2564 1497 2595 1503
rect 980 1477 1027 1483
rect 1044 1477 1084 1483
rect 2404 1477 2444 1483
rect 452 1457 892 1463
rect 900 1457 1196 1463
rect 1636 1457 1788 1463
rect 1796 1457 1804 1463
rect 1828 1457 1948 1463
rect 1812 1437 2076 1443
rect 2084 1437 2188 1443
rect 2196 1437 2236 1443
rect 212 1417 220 1423
rect 228 1417 412 1423
rect 420 1417 492 1423
rect 500 1417 876 1423
rect 884 1417 1260 1423
rect 1620 1417 1660 1423
rect 2052 1417 2492 1423
rect 1858 1414 1918 1416
rect 1858 1406 1859 1414
rect 1868 1406 1869 1414
rect 1907 1406 1908 1414
rect 1917 1406 1918 1414
rect 1858 1404 1918 1406
rect 180 1397 188 1403
rect 2116 1397 2236 1403
rect 580 1377 732 1383
rect 1652 1377 2252 1383
rect 2260 1377 2300 1383
rect 52 1357 108 1363
rect 404 1357 892 1363
rect 900 1357 924 1363
rect 932 1357 1276 1363
rect 1284 1357 1356 1363
rect 1572 1357 1676 1363
rect 2356 1357 2428 1363
rect -35 1337 12 1343
rect 724 1337 924 1343
rect 1108 1337 1388 1343
rect 1492 1337 1564 1343
rect 1604 1337 1612 1343
rect 1716 1337 1772 1343
rect 2164 1337 2204 1343
rect 212 1317 268 1323
rect 484 1317 492 1323
rect 500 1317 812 1323
rect 932 1317 1068 1323
rect 1972 1317 2284 1323
rect 2452 1317 2508 1323
rect -35 1297 60 1303
rect 1012 1297 1068 1303
rect 2100 1297 2156 1303
rect 2308 1297 2364 1303
rect 2228 1277 2412 1283
rect 2420 1277 2444 1283
rect 2468 1277 2508 1283
rect 2020 1257 2124 1263
rect 2132 1257 2172 1263
rect 2276 1257 2380 1263
rect 2404 1257 2444 1263
rect 1236 1237 1276 1243
rect 340 1217 364 1223
rect 1444 1217 1804 1223
rect 642 1214 702 1216
rect 642 1206 643 1214
rect 652 1206 653 1214
rect 691 1206 692 1214
rect 701 1206 702 1214
rect 642 1204 702 1206
rect 308 1197 556 1203
rect 2340 1197 2380 1203
rect 2388 1197 2492 1203
rect 1012 1177 1164 1183
rect 1172 1177 1196 1183
rect 1204 1177 1740 1183
rect 1748 1177 1980 1183
rect 1988 1177 2060 1183
rect 2068 1177 2092 1183
rect 1316 1157 1580 1163
rect 1588 1157 1628 1163
rect 1588 1137 1612 1143
rect 1956 1137 2108 1143
rect 1124 1117 1132 1123
rect 1140 1117 1292 1123
rect 1300 1117 1692 1123
rect 852 1097 892 1103
rect 900 1097 956 1103
rect 1060 1097 1148 1103
rect 1156 1097 1516 1103
rect 1924 1097 1964 1103
rect 2100 1097 2412 1103
rect 196 1077 220 1083
rect 628 1077 908 1083
rect 948 1077 988 1083
rect 1284 1077 1308 1083
rect 1524 1077 1548 1083
rect 1796 1077 1852 1083
rect 1860 1077 2028 1083
rect 2180 1077 2380 1083
rect 909 1063 915 1076
rect 909 1057 972 1063
rect 1108 1057 1244 1063
rect 1316 1057 1564 1063
rect 1572 1057 1676 1063
rect 1684 1057 1772 1063
rect 1780 1057 1804 1063
rect 1124 1037 1324 1043
rect 1476 1037 2012 1043
rect 2020 1037 2076 1043
rect 2084 1037 2172 1043
rect 468 1017 492 1023
rect 1858 1014 1918 1016
rect 1858 1006 1859 1014
rect 1868 1006 1869 1014
rect 1907 1006 1908 1014
rect 1917 1006 1918 1014
rect 1858 1004 1918 1006
rect 100 997 236 1003
rect 244 997 364 1003
rect 372 997 684 1003
rect 692 997 876 1003
rect 1380 997 1468 1003
rect 1540 997 1548 1003
rect 180 977 188 983
rect 196 977 524 983
rect 52 957 108 963
rect 260 957 268 963
rect 276 957 444 963
rect 2212 957 2300 963
rect -35 937 12 943
rect 212 937 220 943
rect 228 937 332 943
rect 356 937 396 943
rect 1652 937 1692 943
rect 1700 937 1740 943
rect 1748 937 1948 943
rect 1956 937 2044 943
rect 2116 937 2124 943
rect 212 917 268 923
rect 308 917 380 923
rect 388 917 428 923
rect 436 917 524 923
rect 532 917 1148 923
rect 1844 917 1964 923
rect 1972 917 2044 923
rect 2420 917 2492 923
rect -35 897 60 903
rect 100 897 364 903
rect 372 897 540 903
rect 548 897 700 903
rect 1460 897 1660 903
rect 1828 897 1964 903
rect 1972 897 1996 903
rect 2004 897 2028 903
rect 2564 897 2595 903
rect 420 877 492 883
rect 1812 877 2428 883
rect 2036 857 2060 863
rect 868 817 940 823
rect 1092 817 1116 823
rect 642 814 702 816
rect 642 806 643 814
rect 652 806 653 814
rect 691 806 692 814
rect 701 806 702 814
rect 642 804 702 806
rect 1668 757 2476 763
rect 420 737 796 743
rect 804 737 924 743
rect 932 737 1132 743
rect 1220 737 1564 743
rect 2148 737 2172 743
rect 2180 737 2252 743
rect 1540 717 1548 723
rect 1716 717 1980 723
rect 1988 717 2012 723
rect 2116 717 2204 723
rect 2212 717 2316 723
rect 324 697 428 703
rect 820 697 844 703
rect 852 697 892 703
rect 900 697 940 703
rect 980 697 1244 703
rect 1508 697 1564 703
rect 1780 697 1820 703
rect 1908 697 2028 703
rect 2100 697 2188 703
rect 2292 697 2460 703
rect 2468 697 2508 703
rect 2564 697 2595 703
rect 196 677 220 683
rect 772 677 876 683
rect 1076 677 1116 683
rect 1524 677 1580 683
rect 1652 677 1708 683
rect 1812 677 1900 683
rect 1924 677 1980 683
rect 1988 677 2044 683
rect 180 657 188 663
rect 388 657 828 663
rect 868 657 924 663
rect 1412 657 1468 663
rect 1476 657 1500 663
rect 1796 657 1932 663
rect 2068 657 2124 663
rect 2196 657 2220 663
rect 2228 657 2252 663
rect 2308 657 2412 663
rect 532 637 780 643
rect 900 637 1116 643
rect 1124 637 1244 643
rect 1252 637 1484 643
rect 1844 637 2060 643
rect 2356 637 2380 643
rect 516 617 556 623
rect 564 617 892 623
rect 2276 617 2444 623
rect 1858 614 1918 616
rect 1858 606 1859 614
rect 1868 606 1869 614
rect 1907 606 1908 614
rect 1917 606 1918 614
rect 1858 604 1918 606
rect 1364 597 1436 603
rect 2468 597 2492 603
rect 2500 597 2508 603
rect 2516 597 2595 603
rect 1556 577 1628 583
rect 2372 577 2396 583
rect -35 557 60 563
rect 68 557 1004 563
rect 1076 557 1100 563
rect 1220 557 1388 563
rect 1396 557 1740 563
rect 1748 557 1836 563
rect 2148 557 2428 563
rect 548 537 620 543
rect 1012 537 1084 543
rect 1716 537 1916 543
rect 2036 537 2092 543
rect 2132 537 2172 543
rect 2180 537 2268 543
rect 2292 537 2332 543
rect 2340 537 2364 543
rect 2436 537 2476 543
rect 2484 537 2595 543
rect 68 517 204 523
rect 308 517 380 523
rect 756 517 844 523
rect 852 517 1020 523
rect 2052 517 2140 523
rect 2148 517 2156 523
rect -35 497 12 503
rect 1988 497 2012 503
rect 2020 497 2204 503
rect 2372 497 2412 503
rect 2589 483 2595 503
rect 2196 477 2595 483
rect 164 457 332 463
rect 340 457 716 463
rect 2388 457 2428 463
rect 356 437 364 443
rect 436 417 476 423
rect 1652 417 1660 423
rect 642 414 702 416
rect 642 406 643 414
rect 652 406 653 414
rect 691 406 692 414
rect 701 406 702 414
rect 642 404 702 406
rect 516 397 572 403
rect 1076 397 1132 403
rect 1396 397 1452 403
rect 660 377 732 383
rect 868 377 924 383
rect 2132 357 2412 363
rect 2420 357 2492 363
rect 2452 337 2492 343
rect -35 317 12 323
rect 724 317 892 323
rect 2132 317 2172 323
rect 100 297 140 303
rect 196 297 204 303
rect 212 297 380 303
rect 884 297 908 303
rect 916 297 1036 303
rect 1268 297 1324 303
rect 1540 297 1628 303
rect 1636 297 1708 303
rect 1940 297 2124 303
rect 2404 297 2556 303
rect 2564 297 2595 303
rect -35 277 92 283
rect 292 277 412 283
rect 1140 277 1148 283
rect 1300 277 1420 283
rect 1428 277 1628 283
rect 2116 277 2204 283
rect 132 257 188 263
rect 2356 257 2460 263
rect 2468 257 2476 263
rect 2484 257 2595 263
rect 1684 237 2140 243
rect 1972 217 2476 223
rect 1858 214 1918 216
rect 1858 206 1859 214
rect 1868 206 1869 214
rect 1907 206 1908 214
rect 1917 206 1918 214
rect 1858 204 1918 206
rect 180 197 220 203
rect 372 197 396 203
rect 404 197 556 203
rect 1556 197 1788 203
rect 2276 197 2412 203
rect 36 177 60 183
rect 548 177 812 183
rect 1812 177 2140 183
rect 2308 177 2332 183
rect 660 157 988 163
rect 1140 157 1452 163
rect 1460 157 1484 163
rect 1780 157 1932 163
rect 1972 157 2012 163
rect 2116 157 2156 163
rect 804 137 860 143
rect 1796 137 2092 143
rect 2100 137 2284 143
rect 2292 137 2316 143
rect 772 117 876 123
rect 1332 117 1356 123
rect 1732 117 1804 123
rect 1956 117 2028 123
rect 2036 117 2172 123
rect 1460 97 1804 103
rect 1924 97 1980 103
rect 2020 97 2156 103
rect 2164 97 2220 103
rect 2244 97 2332 103
rect 2340 97 2380 103
rect 2388 97 2428 103
rect 2564 97 2595 103
rect 2212 77 2252 83
rect 2180 57 2284 63
rect 2148 37 2268 43
rect 642 14 702 16
rect 642 6 643 14
rect 652 6 653 14
rect 691 6 692 14
rect 701 6 702 14
rect 642 4 702 6
<< m4contact >>
rect 364 1816 372 1824
rect 1860 1806 1867 1814
rect 1867 1806 1868 1814
rect 1872 1806 1877 1814
rect 1877 1806 1879 1814
rect 1879 1806 1880 1814
rect 1884 1806 1887 1814
rect 1887 1806 1889 1814
rect 1889 1806 1892 1814
rect 1896 1806 1897 1814
rect 1897 1806 1899 1814
rect 1899 1806 1904 1814
rect 1908 1806 1909 1814
rect 1909 1806 1916 1814
rect 204 1676 212 1684
rect 364 1636 372 1644
rect 1580 1636 1588 1644
rect 644 1606 651 1614
rect 651 1606 652 1614
rect 656 1606 661 1614
rect 661 1606 663 1614
rect 663 1606 664 1614
rect 668 1606 671 1614
rect 671 1606 673 1614
rect 673 1606 676 1614
rect 680 1606 681 1614
rect 681 1606 683 1614
rect 683 1606 688 1614
rect 692 1606 693 1614
rect 693 1606 700 1614
rect 1612 1596 1620 1604
rect 2508 1596 2516 1604
rect 2444 1476 2452 1484
rect 204 1416 212 1424
rect 1860 1406 1867 1414
rect 1867 1406 1868 1414
rect 1872 1406 1877 1414
rect 1877 1406 1879 1414
rect 1879 1406 1880 1414
rect 1884 1406 1887 1414
rect 1887 1406 1889 1414
rect 1889 1406 1892 1414
rect 1896 1406 1897 1414
rect 1897 1406 1899 1414
rect 1899 1406 1904 1414
rect 1908 1406 1909 1414
rect 1909 1406 1916 1414
rect 172 1396 180 1404
rect 1612 1336 1620 1344
rect 2156 1336 2164 1344
rect 268 1316 276 1324
rect 2508 1316 2516 1324
rect 2444 1276 2452 1284
rect 644 1206 651 1214
rect 651 1206 652 1214
rect 656 1206 661 1214
rect 661 1206 663 1214
rect 663 1206 664 1214
rect 668 1206 671 1214
rect 671 1206 673 1214
rect 673 1206 676 1214
rect 680 1206 681 1214
rect 681 1206 683 1214
rect 683 1206 688 1214
rect 692 1206 693 1214
rect 693 1206 700 1214
rect 2380 1196 2388 1204
rect 1580 1156 1588 1164
rect 2028 1056 2036 1064
rect 2156 1016 2164 1024
rect 1860 1006 1867 1014
rect 1867 1006 1868 1014
rect 1872 1006 1877 1014
rect 1877 1006 1879 1014
rect 1879 1006 1880 1014
rect 1884 1006 1887 1014
rect 1887 1006 1889 1014
rect 1889 1006 1892 1014
rect 1896 1006 1897 1014
rect 1897 1006 1899 1014
rect 1899 1006 1904 1014
rect 1908 1006 1909 1014
rect 1909 1006 1916 1014
rect 1548 996 1556 1004
rect 172 976 180 984
rect 268 956 276 964
rect 204 936 212 944
rect 2124 936 2132 944
rect 2028 856 2036 864
rect 644 806 651 814
rect 651 806 652 814
rect 656 806 661 814
rect 661 806 663 814
rect 663 806 664 814
rect 668 806 671 814
rect 671 806 673 814
rect 673 806 676 814
rect 680 806 681 814
rect 681 806 683 814
rect 683 806 688 814
rect 692 806 693 814
rect 693 806 700 814
rect 1548 716 1556 724
rect 1644 696 1652 704
rect 172 656 180 664
rect 1860 606 1867 614
rect 1867 606 1868 614
rect 1872 606 1877 614
rect 1877 606 1879 614
rect 1879 606 1880 614
rect 1884 606 1887 614
rect 1887 606 1889 614
rect 1889 606 1892 614
rect 1896 606 1897 614
rect 1897 606 1899 614
rect 1899 606 1904 614
rect 1908 606 1909 614
rect 1909 606 1916 614
rect 2380 456 2388 464
rect 364 436 372 444
rect 1644 416 1652 424
rect 644 406 651 414
rect 651 406 652 414
rect 656 406 661 414
rect 661 406 663 414
rect 663 406 664 414
rect 668 406 671 414
rect 671 406 673 414
rect 673 406 676 414
rect 680 406 681 414
rect 681 406 683 414
rect 683 406 688 414
rect 692 406 693 414
rect 693 406 700 414
rect 1132 396 1140 404
rect 2124 356 2132 364
rect 1132 276 1140 284
rect 1860 206 1867 214
rect 1867 206 1868 214
rect 1872 206 1877 214
rect 1877 206 1879 214
rect 1879 206 1880 214
rect 1884 206 1887 214
rect 1887 206 1889 214
rect 1889 206 1892 214
rect 1896 206 1897 214
rect 1897 206 1899 214
rect 1899 206 1904 214
rect 1908 206 1909 214
rect 1909 206 1916 214
rect 364 196 372 204
rect 644 6 651 14
rect 651 6 652 14
rect 656 6 661 14
rect 661 6 663 14
rect 663 6 664 14
rect 668 6 671 14
rect 671 6 673 14
rect 673 6 676 14
rect 680 6 681 14
rect 681 6 683 14
rect 683 6 688 14
rect 692 6 693 14
rect 693 6 700 14
<< metal4 >>
rect 362 1824 374 1826
rect 362 1816 364 1824
rect 372 1816 374 1824
rect 202 1684 214 1686
rect 202 1676 204 1684
rect 212 1676 214 1684
rect 202 1424 214 1676
rect 362 1644 374 1816
rect 362 1636 364 1644
rect 372 1636 374 1644
rect 362 1634 374 1636
rect 202 1416 204 1424
rect 212 1416 214 1424
rect 170 1404 182 1406
rect 170 1396 172 1404
rect 180 1396 182 1404
rect 170 984 182 1396
rect 170 976 172 984
rect 180 976 182 984
rect 170 664 182 976
rect 202 944 214 1416
rect 640 1614 704 1816
rect 1856 1814 1920 1816
rect 1856 1806 1860 1814
rect 1868 1806 1872 1814
rect 1880 1806 1884 1814
rect 1892 1806 1896 1814
rect 1904 1806 1908 1814
rect 1916 1806 1920 1814
rect 640 1606 644 1614
rect 652 1606 656 1614
rect 664 1606 668 1614
rect 676 1606 680 1614
rect 688 1606 692 1614
rect 700 1606 704 1614
rect 266 1324 278 1326
rect 266 1316 268 1324
rect 276 1316 278 1324
rect 266 964 278 1316
rect 266 956 268 964
rect 276 956 278 964
rect 266 954 278 956
rect 640 1214 704 1606
rect 640 1206 644 1214
rect 652 1206 656 1214
rect 664 1206 668 1214
rect 676 1206 680 1214
rect 688 1206 692 1214
rect 700 1206 704 1214
rect 202 936 204 944
rect 212 936 214 944
rect 202 934 214 936
rect 170 656 172 664
rect 180 656 182 664
rect 170 654 182 656
rect 640 814 704 1206
rect 1578 1644 1590 1646
rect 1578 1636 1580 1644
rect 1588 1636 1590 1644
rect 1578 1164 1590 1636
rect 1610 1604 1622 1606
rect 1610 1596 1612 1604
rect 1620 1596 1622 1604
rect 1610 1344 1622 1596
rect 1610 1336 1612 1344
rect 1620 1336 1622 1344
rect 1610 1334 1622 1336
rect 1856 1414 1920 1806
rect 2506 1604 2518 1606
rect 2506 1596 2508 1604
rect 2516 1596 2518 1604
rect 1856 1406 1860 1414
rect 1868 1406 1872 1414
rect 1880 1406 1884 1414
rect 1892 1406 1896 1414
rect 1904 1406 1908 1414
rect 1916 1406 1920 1414
rect 1578 1156 1580 1164
rect 1588 1156 1590 1164
rect 1578 1154 1590 1156
rect 1856 1014 1920 1406
rect 2442 1484 2454 1486
rect 2442 1476 2444 1484
rect 2452 1476 2454 1484
rect 2154 1344 2166 1346
rect 2154 1336 2156 1344
rect 2164 1336 2166 1344
rect 1856 1006 1860 1014
rect 1868 1006 1872 1014
rect 1880 1006 1884 1014
rect 1892 1006 1896 1014
rect 1904 1006 1908 1014
rect 1916 1006 1920 1014
rect 640 806 644 814
rect 652 806 656 814
rect 664 806 668 814
rect 676 806 680 814
rect 688 806 692 814
rect 700 806 704 814
rect 362 444 374 446
rect 362 436 364 444
rect 372 436 374 444
rect 362 204 374 436
rect 362 196 364 204
rect 372 196 374 204
rect 362 194 374 196
rect 640 414 704 806
rect 1546 1004 1558 1006
rect 1546 996 1548 1004
rect 1556 996 1558 1004
rect 1546 724 1558 996
rect 1546 716 1548 724
rect 1556 716 1558 724
rect 1546 714 1558 716
rect 1642 704 1654 706
rect 1642 696 1644 704
rect 1652 696 1654 704
rect 1642 424 1654 696
rect 1642 416 1644 424
rect 1652 416 1654 424
rect 1642 414 1654 416
rect 1856 614 1920 1006
rect 2026 1064 2038 1066
rect 2026 1056 2028 1064
rect 2036 1056 2038 1064
rect 2026 864 2038 1056
rect 2154 1024 2166 1336
rect 2442 1284 2454 1476
rect 2506 1324 2518 1596
rect 2506 1316 2508 1324
rect 2516 1316 2518 1324
rect 2506 1314 2518 1316
rect 2442 1276 2444 1284
rect 2452 1276 2454 1284
rect 2442 1274 2454 1276
rect 2154 1016 2156 1024
rect 2164 1016 2166 1024
rect 2154 1014 2166 1016
rect 2378 1204 2390 1206
rect 2378 1196 2380 1204
rect 2388 1196 2390 1204
rect 2026 856 2028 864
rect 2036 856 2038 864
rect 2026 854 2038 856
rect 2122 944 2134 946
rect 2122 936 2124 944
rect 2132 936 2134 944
rect 1856 606 1860 614
rect 1868 606 1872 614
rect 1880 606 1884 614
rect 1892 606 1896 614
rect 1904 606 1908 614
rect 1916 606 1920 614
rect 640 406 644 414
rect 652 406 656 414
rect 664 406 668 414
rect 676 406 680 414
rect 688 406 692 414
rect 700 406 704 414
rect 640 14 704 406
rect 1130 404 1142 406
rect 1130 396 1132 404
rect 1140 396 1142 404
rect 1130 284 1142 396
rect 1130 276 1132 284
rect 1140 276 1142 284
rect 1130 274 1142 276
rect 640 6 644 14
rect 652 6 656 14
rect 664 6 668 14
rect 676 6 680 14
rect 688 6 692 14
rect 700 6 704 14
rect 640 -10 704 6
rect 1856 214 1920 606
rect 2122 364 2134 936
rect 2378 464 2390 1196
rect 2378 456 2380 464
rect 2388 456 2390 464
rect 2378 454 2390 456
rect 2122 356 2124 364
rect 2132 356 2134 364
rect 2122 354 2134 356
rect 1856 206 1860 214
rect 1868 206 1872 214
rect 1880 206 1884 214
rect 1892 206 1896 214
rect 1904 206 1908 214
rect 1916 206 1920 214
rect 1856 -10 1920 206
use BUFX2  _265_
timestamp 1593098107
transform -1 0 56 0 -1 1810
box -4 -6 52 206
use INVX1  _150_
timestamp 1593098107
transform 1 0 56 0 -1 1810
box -4 -6 36 206
use MUX2X1  _152_
timestamp 1593098107
transform -1 0 184 0 -1 1810
box -4 -6 100 206
use DFFSR  _298_
timestamp 1593098107
transform 1 0 184 0 -1 1810
box -4 -6 356 206
use BUFX2  _258_
timestamp 1593098107
transform 1 0 536 0 -1 1810
box -4 -6 52 206
use BUFX2  _273_
timestamp 1593098107
transform 1 0 584 0 -1 1810
box -4 -6 52 206
use FILL  SFILL6320x16100
timestamp 1593098107
transform -1 0 648 0 -1 1810
box -4 -6 20 206
use FILL  SFILL6480x16100
timestamp 1593098107
transform -1 0 664 0 -1 1810
box -4 -6 20 206
use FILL  SFILL6640x16100
timestamp 1593098107
transform -1 0 680 0 -1 1810
box -4 -6 20 206
use FILL  SFILL6800x16100
timestamp 1593098107
transform -1 0 696 0 -1 1810
box -4 -6 20 206
use BUFX2  _259_
timestamp 1593098107
transform -1 0 744 0 -1 1810
box -4 -6 52 206
use DFFSR  _299_
timestamp 1593098107
transform -1 0 1096 0 -1 1810
box -4 -6 356 206
use INVX8  _247_
timestamp 1593098107
transform 1 0 1096 0 -1 1810
box -4 -6 84 206
use DFFSR  _278_
timestamp 1593098107
transform 1 0 1176 0 -1 1810
box -4 -6 356 206
use BUFX2  _256_
timestamp 1593098107
transform -1 0 1576 0 -1 1810
box -4 -6 52 206
use INVX1  _176_
timestamp 1593098107
transform 1 0 1576 0 -1 1810
box -4 -6 36 206
use DFFSR  _276_
timestamp 1593098107
transform -1 0 1960 0 -1 1810
box -4 -6 356 206
use FILL  SFILL19600x16100
timestamp 1593098107
transform -1 0 1976 0 -1 1810
box -4 -6 20 206
use FILL  SFILL19760x16100
timestamp 1593098107
transform -1 0 1992 0 -1 1810
box -4 -6 20 206
use FILL  SFILL19920x16100
timestamp 1593098107
transform -1 0 2008 0 -1 1810
box -4 -6 20 206
use FILL  SFILL20080x16100
timestamp 1593098107
transform -1 0 2024 0 -1 1810
box -4 -6 20 206
use BUFX2  _255_
timestamp 1593098107
transform 1 0 2024 0 -1 1810
box -4 -6 52 206
use DFFSR  _287_
timestamp 1593098107
transform 1 0 2072 0 -1 1810
box -4 -6 356 206
use OAI21X1  _237_
timestamp 1593098107
transform 1 0 2424 0 -1 1810
box -4 -6 68 206
use INVX1  _236_
timestamp 1593098107
transform -1 0 2520 0 -1 1810
box -4 -6 36 206
use FILL  FILL23920x16100
timestamp 1593098107
transform -1 0 2536 0 -1 1810
box -4 -6 20 206
use FILL  FILL24080x16100
timestamp 1593098107
transform -1 0 2552 0 -1 1810
box -4 -6 20 206
use DFFSR  _305_
timestamp 1593098107
transform -1 0 360 0 1 1410
box -4 -6 356 206
use BUFX2  _266_
timestamp 1593098107
transform -1 0 408 0 1 1410
box -4 -6 52 206
use NOR2X1  _130_
timestamp 1593098107
transform -1 0 456 0 1 1410
box -4 -6 52 206
use AOI21X1  _131_
timestamp 1593098107
transform -1 0 520 0 1 1410
box -4 -6 68 206
use INVX1  _127_
timestamp 1593098107
transform -1 0 552 0 1 1410
box -4 -6 36 206
use INVX1  _151_
timestamp 1593098107
transform -1 0 584 0 1 1410
box -4 -6 36 206
use BUFX2  _272_
timestamp 1593098107
transform 1 0 584 0 1 1410
box -4 -6 52 206
use FILL  SFILL6320x14100
timestamp 1593098107
transform 1 0 632 0 1 1410
box -4 -6 20 206
use FILL  SFILL6480x14100
timestamp 1593098107
transform 1 0 648 0 1 1410
box -4 -6 20 206
use FILL  SFILL6640x14100
timestamp 1593098107
transform 1 0 664 0 1 1410
box -4 -6 20 206
use FILL  SFILL6800x14100
timestamp 1593098107
transform 1 0 680 0 1 1410
box -4 -6 20 206
use AOI21X1  _173_
timestamp 1593098107
transform -1 0 760 0 1 1410
box -4 -6 68 206
use INVX1  _132_
timestamp 1593098107
transform 1 0 760 0 1 1410
box -4 -6 36 206
use MUX2X1  _134_
timestamp 1593098107
transform -1 0 888 0 1 1410
box -4 -6 100 206
use OAI21X1  _174_
timestamp 1593098107
transform 1 0 888 0 1 1410
box -4 -6 68 206
use AOI21X1  _175_
timestamp 1593098107
transform -1 0 1016 0 1 1410
box -4 -6 68 206
use INVX1  _133_
timestamp 1593098107
transform -1 0 1048 0 1 1410
box -4 -6 36 206
use BUFX2  _267_
timestamp 1593098107
transform -1 0 1096 0 1 1410
box -4 -6 52 206
use DFFSR  _290_
timestamp 1593098107
transform -1 0 1448 0 1 1410
box -4 -6 356 206
use DFFSR  _306_
timestamp 1593098107
transform -1 0 1800 0 1 1410
box -4 -6 356 206
use INVX1  _246_
timestamp 1593098107
transform -1 0 1832 0 1 1410
box -4 -6 36 206
use FILL  SFILL18320x14100
timestamp 1593098107
transform 1 0 1832 0 1 1410
box -4 -6 20 206
use FILL  SFILL18480x14100
timestamp 1593098107
transform 1 0 1848 0 1 1410
box -4 -6 20 206
use FILL  SFILL18640x14100
timestamp 1593098107
transform 1 0 1864 0 1 1410
box -4 -6 20 206
use FILL  SFILL18800x14100
timestamp 1593098107
transform 1 0 1880 0 1 1410
box -4 -6 20 206
use DFFSR  _288_
timestamp 1593098107
transform -1 0 2248 0 1 1410
box -4 -6 356 206
use OAI21X1  _235_
timestamp 1593098107
transform 1 0 2248 0 1 1410
box -4 -6 68 206
use INVX1  _227_
timestamp 1593098107
transform 1 0 2312 0 1 1410
box -4 -6 36 206
use OAI21X1  _228_
timestamp 1593098107
transform -1 0 2408 0 1 1410
box -4 -6 68 206
use INVX1  _224_
timestamp 1593098107
transform -1 0 2440 0 1 1410
box -4 -6 36 206
use BUFX2  _254_
timestamp 1593098107
transform 1 0 2440 0 1 1410
box -4 -6 52 206
use BUFX2  _248_
timestamp 1593098107
transform 1 0 2488 0 1 1410
box -4 -6 52 206
use FILL  FILL24080x14100
timestamp 1593098107
transform 1 0 2536 0 1 1410
box -4 -6 20 206
use BUFX2  _263_
timestamp 1593098107
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use BUFX2  _271_
timestamp 1593098107
transform -1 0 104 0 -1 1410
box -4 -6 52 206
use INVX1  _144_
timestamp 1593098107
transform 1 0 104 0 -1 1410
box -4 -6 36 206
use MUX2X1  _146_
timestamp 1593098107
transform -1 0 232 0 -1 1410
box -4 -6 100 206
use DFFSR  _295_
timestamp 1593098107
transform 1 0 232 0 -1 1410
box -4 -6 356 206
use OAI21X1  _172_
timestamp 1593098107
transform 1 0 584 0 -1 1410
box -4 -6 68 206
use FILL  SFILL6480x12100
timestamp 1593098107
transform -1 0 664 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6640x12100
timestamp 1593098107
transform -1 0 680 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6800x12100
timestamp 1593098107
transform -1 0 696 0 -1 1410
box -4 -6 20 206
use FILL  SFILL6960x12100
timestamp 1593098107
transform -1 0 712 0 -1 1410
box -4 -6 20 206
use DFFSR  _296_
timestamp 1593098107
transform -1 0 1064 0 -1 1410
box -4 -6 356 206
use NOR2X1  _161_
timestamp 1593098107
transform -1 0 1112 0 -1 1410
box -4 -6 52 206
use OAI21X1  _160_
timestamp 1593098107
transform -1 0 1176 0 -1 1410
box -4 -6 68 206
use DFFSR  _289_
timestamp 1593098107
transform -1 0 1528 0 -1 1410
box -4 -6 356 206
use BUFX2  BUFX2_insert12
timestamp 1593098107
transform 1 0 1528 0 -1 1410
box -4 -6 52 206
use AOI21X1  _179_
timestamp 1593098107
transform 1 0 1576 0 -1 1410
box -4 -6 68 206
use DFFSR  _277_
timestamp 1593098107
transform 1 0 1640 0 -1 1410
box -4 -6 356 206
use FILL  SFILL19920x12100
timestamp 1593098107
transform -1 0 2008 0 -1 1410
box -4 -6 20 206
use FILL  SFILL20080x12100
timestamp 1593098107
transform -1 0 2024 0 -1 1410
box -4 -6 20 206
use FILL  SFILL20240x12100
timestamp 1593098107
transform -1 0 2040 0 -1 1410
box -4 -6 20 206
use FILL  SFILL20400x12100
timestamp 1593098107
transform -1 0 2056 0 -1 1410
box -4 -6 20 206
use INVX1  _240_
timestamp 1593098107
transform 1 0 2056 0 -1 1410
box -4 -6 36 206
use NAND3X1  _241_
timestamp 1593098107
transform 1 0 2088 0 -1 1410
box -4 -6 68 206
use AOI22X1  _234_
timestamp 1593098107
transform 1 0 2152 0 -1 1410
box -4 -6 84 206
use AND2X2  _244_
timestamp 1593098107
transform -1 0 2296 0 -1 1410
box -4 -6 68 206
use OAI21X1  _226_
timestamp 1593098107
transform -1 0 2360 0 -1 1410
box -4 -6 68 206
use NAND3X1  _239_
timestamp 1593098107
transform 1 0 2360 0 -1 1410
box -4 -6 68 206
use NAND3X1  _238_
timestamp 1593098107
transform 1 0 2424 0 -1 1410
box -4 -6 68 206
use INVX1  _225_
timestamp 1593098107
transform 1 0 2488 0 -1 1410
box -4 -6 36 206
use FILL  FILL23920x12100
timestamp 1593098107
transform -1 0 2536 0 -1 1410
box -4 -6 20 206
use FILL  FILL24080x12100
timestamp 1593098107
transform -1 0 2552 0 -1 1410
box -4 -6 20 206
use DFFSR  _303_
timestamp 1593098107
transform -1 0 360 0 1 1010
box -4 -6 356 206
use DFFSR  _294_
timestamp 1593098107
transform 1 0 360 0 1 1010
box -4 -6 356 206
use FILL  SFILL7120x10100
timestamp 1593098107
transform 1 0 712 0 1 1010
box -4 -6 20 206
use FILL  SFILL7280x10100
timestamp 1593098107
transform 1 0 728 0 1 1010
box -4 -6 20 206
use FILL  SFILL7440x10100
timestamp 1593098107
transform 1 0 744 0 1 1010
box -4 -6 20 206
use FILL  SFILL7600x10100
timestamp 1593098107
transform 1 0 760 0 1 1010
box -4 -6 20 206
use XNOR2X1  _156_
timestamp 1593098107
transform -1 0 888 0 1 1010
box -4 -6 116 206
use AOI21X1  _159_
timestamp 1593098107
transform 1 0 888 0 1 1010
box -4 -6 68 206
use OAI21X1  _158_
timestamp 1593098107
transform 1 0 952 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert9
timestamp 1593098107
transform -1 0 1064 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert7
timestamp 1593098107
transform -1 0 1112 0 1 1010
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert0
timestamp 1593098107
transform 1 0 1112 0 1 1010
box -4 -6 148 206
use NAND3X1  _129_
timestamp 1593098107
transform -1 0 1320 0 1 1010
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert1
timestamp 1593098107
transform 1 0 1320 0 1 1010
box -4 -6 148 206
use BUFX2  BUFX2_insert13
timestamp 1593098107
transform -1 0 1512 0 1 1010
box -4 -6 52 206
use INVX1  _123_
timestamp 1593098107
transform 1 0 1512 0 1 1010
box -4 -6 36 206
use NAND3X1  _178_
timestamp 1593098107
transform 1 0 1544 0 1 1010
box -4 -6 68 206
use INVX1  _177_
timestamp 1593098107
transform -1 0 1640 0 1 1010
box -4 -6 36 206
use INVX4  _115_
timestamp 1593098107
transform 1 0 1640 0 1 1010
box -4 -6 52 206
use NAND2X1  _121_
timestamp 1593098107
transform 1 0 1688 0 1 1010
box -4 -6 52 206
use OAI21X1  _120_
timestamp 1593098107
transform -1 0 1800 0 1 1010
box -4 -6 68 206
use OAI21X1  _242_
timestamp 1593098107
transform 1 0 1800 0 1 1010
box -4 -6 68 206
use FILL  SFILL18640x10100
timestamp 1593098107
transform 1 0 1864 0 1 1010
box -4 -6 20 206
use FILL  SFILL18800x10100
timestamp 1593098107
transform 1 0 1880 0 1 1010
box -4 -6 20 206
use FILL  SFILL18960x10100
timestamp 1593098107
transform 1 0 1896 0 1 1010
box -4 -6 20 206
use FILL  SFILL19120x10100
timestamp 1593098107
transform 1 0 1912 0 1 1010
box -4 -6 20 206
use NAND3X1  _243_
timestamp 1593098107
transform -1 0 1992 0 1 1010
box -4 -6 68 206
use NOR2X1  _232_
timestamp 1593098107
transform -1 0 2040 0 1 1010
box -4 -6 52 206
use DFFSR  _286_
timestamp 1593098107
transform 1 0 2040 0 1 1010
box -4 -6 356 206
use NOR3X1  _118_
timestamp 1593098107
transform 1 0 2392 0 1 1010
box -4 -6 132 206
use FILL  FILL23920x10100
timestamp 1593098107
transform 1 0 2520 0 1 1010
box -4 -6 20 206
use FILL  FILL24080x10100
timestamp 1593098107
transform 1 0 2536 0 1 1010
box -4 -6 20 206
use BUFX2  _264_
timestamp 1593098107
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use BUFX2  _270_
timestamp 1593098107
transform -1 0 104 0 -1 1010
box -4 -6 52 206
use INVX1  _147_
timestamp 1593098107
transform 1 0 104 0 -1 1010
box -4 -6 36 206
use MUX2X1  _149_
timestamp 1593098107
transform -1 0 232 0 -1 1010
box -4 -6 100 206
use INVX1  _145_
timestamp 1593098107
transform 1 0 232 0 -1 1010
box -4 -6 36 206
use INVX1  _148_
timestamp 1593098107
transform -1 0 296 0 -1 1010
box -4 -6 36 206
use AOI21X1  _171_
timestamp 1593098107
transform 1 0 296 0 -1 1010
box -4 -6 68 206
use OAI21X1  _170_
timestamp 1593098107
transform 1 0 360 0 -1 1010
box -4 -6 68 206
use AOI21X1  _169_
timestamp 1593098107
transform 1 0 424 0 -1 1010
box -4 -6 68 206
use OAI21X1  _168_
timestamp 1593098107
transform -1 0 552 0 -1 1010
box -4 -6 68 206
use XNOR2X1  _157_
timestamp 1593098107
transform -1 0 664 0 -1 1010
box -4 -6 116 206
use FILL  SFILL6640x8100
timestamp 1593098107
transform -1 0 680 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6800x8100
timestamp 1593098107
transform -1 0 696 0 -1 1010
box -4 -6 20 206
use FILL  SFILL6960x8100
timestamp 1593098107
transform -1 0 712 0 -1 1010
box -4 -6 20 206
use FILL  SFILL7120x8100
timestamp 1593098107
transform -1 0 728 0 -1 1010
box -4 -6 20 206
use DFFSR  _293_
timestamp 1593098107
transform -1 0 1080 0 -1 1010
box -4 -6 356 206
use OAI21X1  _162_
timestamp 1593098107
transform 1 0 1080 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert8
timestamp 1593098107
transform -1 0 1192 0 -1 1010
box -4 -6 52 206
use INVX8  _128_
timestamp 1593098107
transform 1 0 1192 0 -1 1010
box -4 -6 84 206
use BUFX2  BUFX2_insert5
timestamp 1593098107
transform 1 0 1272 0 -1 1010
box -4 -6 52 206
use DFFSR  _281_
timestamp 1593098107
transform 1 0 1320 0 -1 1010
box -4 -6 356 206
use AND2X2  _181_
timestamp 1593098107
transform 1 0 1672 0 -1 1010
box -4 -6 68 206
use NOR2X1  _182_
timestamp 1593098107
transform 1 0 1736 0 -1 1010
box -4 -6 52 206
use NAND3X1  _119_
timestamp 1593098107
transform -1 0 1848 0 -1 1010
box -4 -6 68 206
use FILL  SFILL18480x8100
timestamp 1593098107
transform -1 0 1864 0 -1 1010
box -4 -6 20 206
use FILL  SFILL18640x8100
timestamp 1593098107
transform -1 0 1880 0 -1 1010
box -4 -6 20 206
use FILL  SFILL18800x8100
timestamp 1593098107
transform -1 0 1896 0 -1 1010
box -4 -6 20 206
use FILL  SFILL18960x8100
timestamp 1593098107
transform -1 0 1912 0 -1 1010
box -4 -6 20 206
use NOR2X1  _117_
timestamp 1593098107
transform 1 0 1912 0 -1 1010
box -4 -6 52 206
use NAND2X1  _229_
timestamp 1593098107
transform 1 0 1960 0 -1 1010
box -4 -6 52 206
use NAND3X1  _204_
timestamp 1593098107
transform -1 0 2072 0 -1 1010
box -4 -6 68 206
use INVX1  _230_
timestamp 1593098107
transform -1 0 2104 0 -1 1010
box -4 -6 36 206
use INVX2  _187_
timestamp 1593098107
transform 1 0 2104 0 -1 1010
box -4 -6 36 206
use DFFSR  _285_
timestamp 1593098107
transform 1 0 2136 0 -1 1010
box -4 -6 356 206
use BUFX2  _253_
timestamp 1593098107
transform 1 0 2488 0 -1 1010
box -4 -6 52 206
use FILL  FILL24080x8100
timestamp 1593098107
transform -1 0 2552 0 -1 1010
box -4 -6 20 206
use DFFSR  _304_
timestamp 1593098107
transform -1 0 360 0 1 610
box -4 -6 356 206
use INVX1  _142_
timestamp 1593098107
transform 1 0 360 0 1 610
box -4 -6 36 206
use DFFSR  _292_
timestamp 1593098107
transform 1 0 392 0 1 610
box -4 -6 356 206
use FILL  SFILL7440x6100
timestamp 1593098107
transform 1 0 744 0 1 610
box -4 -6 20 206
use FILL  SFILL7600x6100
timestamp 1593098107
transform 1 0 760 0 1 610
box -4 -6 20 206
use FILL  SFILL7760x6100
timestamp 1593098107
transform 1 0 776 0 1 610
box -4 -6 20 206
use FILL  SFILL7920x6100
timestamp 1593098107
transform 1 0 792 0 1 610
box -4 -6 20 206
use AOI21X1  _167_
timestamp 1593098107
transform 1 0 808 0 1 610
box -4 -6 68 206
use OAI21X1  _166_
timestamp 1593098107
transform 1 0 872 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert6
timestamp 1593098107
transform -1 0 984 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert10
timestamp 1593098107
transform -1 0 1032 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert11
timestamp 1593098107
transform 1 0 1032 0 1 610
box -4 -6 52 206
use DFFSR  _275_
timestamp 1593098107
transform 1 0 1080 0 1 610
box -4 -6 356 206
use AND2X2  _245_
timestamp 1593098107
transform -1 0 1496 0 1 610
box -4 -6 68 206
use INVX1  _122_
timestamp 1593098107
transform 1 0 1496 0 1 610
box -4 -6 36 206
use OAI21X1  _126_
timestamp 1593098107
transform -1 0 1592 0 1 610
box -4 -6 68 206
use NOR2X1  _125_
timestamp 1593098107
transform 1 0 1592 0 1 610
box -4 -6 52 206
use OAI21X1  _184_
timestamp 1593098107
transform 1 0 1640 0 1 610
box -4 -6 68 206
use OAI21X1  _183_
timestamp 1593098107
transform -1 0 1768 0 1 610
box -4 -6 68 206
use NAND2X1  _190_
timestamp 1593098107
transform -1 0 1816 0 1 610
box -4 -6 52 206
use NOR2X1  _192_
timestamp 1593098107
transform -1 0 1864 0 1 610
box -4 -6 52 206
use FILL  SFILL18640x6100
timestamp 1593098107
transform 1 0 1864 0 1 610
box -4 -6 20 206
use FILL  SFILL18800x6100
timestamp 1593098107
transform 1 0 1880 0 1 610
box -4 -6 20 206
use FILL  SFILL18960x6100
timestamp 1593098107
transform 1 0 1896 0 1 610
box -4 -6 20 206
use FILL  SFILL19120x6100
timestamp 1593098107
transform 1 0 1912 0 1 610
box -4 -6 20 206
use INVX1  _191_
timestamp 1593098107
transform 1 0 1928 0 1 610
box -4 -6 36 206
use OAI21X1  _193_
timestamp 1593098107
transform 1 0 1960 0 1 610
box -4 -6 68 206
use INVX1  _189_
timestamp 1593098107
transform -1 0 2056 0 1 610
box -4 -6 36 206
use NAND3X1  _231_
timestamp 1593098107
transform -1 0 2120 0 1 610
box -4 -6 68 206
use INVX1  _211_
timestamp 1593098107
transform 1 0 2120 0 1 610
box -4 -6 36 206
use NAND3X1  _233_
timestamp 1593098107
transform -1 0 2216 0 1 610
box -4 -6 68 206
use NOR2X1  _212_
timestamp 1593098107
transform 1 0 2216 0 1 610
box -4 -6 52 206
use INVX1  _210_
timestamp 1593098107
transform -1 0 2296 0 1 610
box -4 -6 36 206
use INVX1  _221_
timestamp 1593098107
transform 1 0 2296 0 1 610
box -4 -6 36 206
use AOI22X1  _223_
timestamp 1593098107
transform 1 0 2328 0 1 610
box -4 -6 84 206
use OAI21X1  _220_
timestamp 1593098107
transform -1 0 2472 0 1 610
box -4 -6 68 206
use INVX1  _180_
timestamp 1593098107
transform -1 0 2504 0 1 610
box -4 -6 36 206
use BUFX2  _252_
timestamp 1593098107
transform 1 0 2504 0 1 610
box -4 -6 52 206
use BUFX2  _262_
timestamp 1593098107
transform -1 0 56 0 -1 610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert4
timestamp 1593098107
transform 1 0 56 0 -1 610
box -4 -6 148 206
use INVX1  _141_
timestamp 1593098107
transform 1 0 200 0 -1 610
box -4 -6 36 206
use MUX2X1  _143_
timestamp 1593098107
transform -1 0 328 0 -1 610
box -4 -6 100 206
use DFFSR  _301_
timestamp 1593098107
transform -1 0 680 0 -1 610
box -4 -6 356 206
use FILL  SFILL6800x4100
timestamp 1593098107
transform -1 0 696 0 -1 610
box -4 -6 20 206
use FILL  SFILL6960x4100
timestamp 1593098107
transform -1 0 712 0 -1 610
box -4 -6 20 206
use FILL  SFILL7120x4100
timestamp 1593098107
transform -1 0 728 0 -1 610
box -4 -6 20 206
use FILL  SFILL7280x4100
timestamp 1593098107
transform -1 0 744 0 -1 610
box -4 -6 20 206
use AOI21X1  _165_
timestamp 1593098107
transform 1 0 744 0 -1 610
box -4 -6 68 206
use OAI21X1  _164_
timestamp 1593098107
transform -1 0 872 0 -1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert2
timestamp 1593098107
transform -1 0 1016 0 -1 610
box -4 -6 148 206
use AOI21X1  _163_
timestamp 1593098107
transform 1 0 1016 0 -1 610
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert3
timestamp 1593098107
transform 1 0 1080 0 -1 610
box -4 -6 148 206
use DFFSR  _274_
timestamp 1593098107
transform 1 0 1224 0 -1 610
box -4 -6 356 206
use DFFSR  _282_
timestamp 1593098107
transform 1 0 1576 0 -1 610
box -4 -6 356 206
use FILL  SFILL19280x4100
timestamp 1593098107
transform -1 0 1944 0 -1 610
box -4 -6 20 206
use FILL  SFILL19440x4100
timestamp 1593098107
transform -1 0 1960 0 -1 610
box -4 -6 20 206
use FILL  SFILL19600x4100
timestamp 1593098107
transform -1 0 1976 0 -1 610
box -4 -6 20 206
use FILL  SFILL19760x4100
timestamp 1593098107
transform -1 0 1992 0 -1 610
box -4 -6 20 206
use NAND2X1  _194_
timestamp 1593098107
transform -1 0 2040 0 -1 610
box -4 -6 52 206
use NOR2X1  _116_
timestamp 1593098107
transform -1 0 2088 0 -1 610
box -4 -6 52 206
use OAI21X1  _188_
timestamp 1593098107
transform -1 0 2152 0 -1 610
box -4 -6 68 206
use BUFX2  _250_
timestamp 1593098107
transform 1 0 2152 0 -1 610
box -4 -6 52 206
use OAI21X1  _214_
timestamp 1593098107
transform -1 0 2264 0 -1 610
box -4 -6 68 206
use NOR2X1  _213_
timestamp 1593098107
transform -1 0 2312 0 -1 610
box -4 -6 52 206
use AOI21X1  _222_
timestamp 1593098107
transform 1 0 2312 0 -1 610
box -4 -6 68 206
use NAND2X1  _219_
timestamp 1593098107
transform 1 0 2376 0 -1 610
box -4 -6 52 206
use NOR2X1  _185_
timestamp 1593098107
transform -1 0 2472 0 -1 610
box -4 -6 52 206
use NAND2X1  _186_
timestamp 1593098107
transform -1 0 2520 0 -1 610
box -4 -6 52 206
use FILL  FILL23920x4100
timestamp 1593098107
transform -1 0 2536 0 -1 610
box -4 -6 20 206
use FILL  FILL24080x4100
timestamp 1593098107
transform -1 0 2552 0 -1 610
box -4 -6 20 206
use BUFX2  _257_
timestamp 1593098107
transform -1 0 56 0 1 210
box -4 -6 52 206
use INVX1  _153_
timestamp 1593098107
transform 1 0 56 0 1 210
box -4 -6 36 206
use NOR2X1  _154_
timestamp 1593098107
transform 1 0 88 0 1 210
box -4 -6 52 206
use AOI21X1  _155_
timestamp 1593098107
transform 1 0 136 0 1 210
box -4 -6 68 206
use DFFSR  _302_
timestamp 1593098107
transform -1 0 552 0 1 210
box -4 -6 356 206
use INVX1  _138_
timestamp 1593098107
transform 1 0 552 0 1 210
box -4 -6 36 206
use MUX2X1  _140_
timestamp 1593098107
transform -1 0 680 0 1 210
box -4 -6 100 206
use FILL  SFILL6800x2100
timestamp 1593098107
transform 1 0 680 0 1 210
box -4 -6 20 206
use FILL  SFILL6960x2100
timestamp 1593098107
transform 1 0 696 0 1 210
box -4 -6 20 206
use FILL  SFILL7120x2100
timestamp 1593098107
transform 1 0 712 0 1 210
box -4 -6 20 206
use FILL  SFILL7280x2100
timestamp 1593098107
transform 1 0 728 0 1 210
box -4 -6 20 206
use INVX1  _139_
timestamp 1593098107
transform -1 0 776 0 1 210
box -4 -6 36 206
use INVX1  _135_
timestamp 1593098107
transform -1 0 808 0 1 210
box -4 -6 36 206
use MUX2X1  _137_
timestamp 1593098107
transform -1 0 904 0 1 210
box -4 -6 100 206
use INVX1  _136_
timestamp 1593098107
transform -1 0 936 0 1 210
box -4 -6 36 206
use DFFSR  _291_
timestamp 1593098107
transform -1 0 1288 0 1 210
box -4 -6 356 206
use DFFSR  _280_
timestamp 1593098107
transform 1 0 1288 0 1 210
box -4 -6 356 206
use INVX1  _124_
timestamp 1593098107
transform 1 0 1640 0 1 210
box -4 -6 36 206
use DFFSR  _284_
timestamp 1593098107
transform 1 0 1672 0 1 210
box -4 -6 356 206
use FILL  SFILL20240x2100
timestamp 1593098107
transform 1 0 2024 0 1 210
box -4 -6 20 206
use FILL  SFILL20400x2100
timestamp 1593098107
transform 1 0 2040 0 1 210
box -4 -6 20 206
use FILL  SFILL20560x2100
timestamp 1593098107
transform 1 0 2056 0 1 210
box -4 -6 20 206
use FILL  SFILL20720x2100
timestamp 1593098107
transform 1 0 2072 0 1 210
box -4 -6 20 206
use OAI21X1  _203_
timestamp 1593098107
transform -1 0 2152 0 1 210
box -4 -6 68 206
use AND2X2  _205_
timestamp 1593098107
transform -1 0 2216 0 1 210
box -4 -6 68 206
use OAI21X1  _215_
timestamp 1593098107
transform -1 0 2280 0 1 210
box -4 -6 68 206
use OAI21X1  _209_
timestamp 1593098107
transform -1 0 2344 0 1 210
box -4 -6 68 206
use OAI21X1  _218_
timestamp 1593098107
transform 1 0 2344 0 1 210
box -4 -6 68 206
use NAND3X1  _217_
timestamp 1593098107
transform 1 0 2408 0 1 210
box -4 -6 68 206
use NOR2X1  _216_
timestamp 1593098107
transform 1 0 2472 0 1 210
box -4 -6 52 206
use FILL  FILL23920x2100
timestamp 1593098107
transform 1 0 2520 0 1 210
box -4 -6 20 206
use FILL  FILL24080x2100
timestamp 1593098107
transform 1 0 2536 0 1 210
box -4 -6 20 206
use DFFSR  _297_
timestamp 1593098107
transform -1 0 360 0 -1 210
box -4 -6 356 206
use BUFX2  _261_
timestamp 1593098107
transform -1 0 408 0 -1 210
box -4 -6 52 206
use DFFSR  _300_
timestamp 1593098107
transform 1 0 408 0 -1 210
box -4 -6 356 206
use FILL  SFILL7600x100
timestamp 1593098107
transform -1 0 776 0 -1 210
box -4 -6 20 206
use FILL  SFILL7760x100
timestamp 1593098107
transform -1 0 792 0 -1 210
box -4 -6 20 206
use FILL  SFILL7920x100
timestamp 1593098107
transform -1 0 808 0 -1 210
box -4 -6 20 206
use FILL  SFILL8080x100
timestamp 1593098107
transform -1 0 824 0 -1 210
box -4 -6 20 206
use BUFX2  _260_
timestamp 1593098107
transform -1 0 872 0 -1 210
box -4 -6 52 206
use BUFX2  _269_
timestamp 1593098107
transform 1 0 872 0 -1 210
box -4 -6 52 206
use BUFX2  _268_
timestamp 1593098107
transform 1 0 920 0 -1 210
box -4 -6 52 206
use DFFSR  _279_
timestamp 1593098107
transform 1 0 968 0 -1 210
box -4 -6 356 206
use DFFSR  _283_
timestamp 1593098107
transform 1 0 1320 0 -1 210
box -4 -6 356 206
use XOR2X1  _197_
timestamp 1593098107
transform -1 0 1784 0 -1 210
box -4 -6 116 206
use OAI21X1  _198_
timestamp 1593098107
transform 1 0 1784 0 -1 210
box -4 -6 68 206
use FILL  SFILL18480x100
timestamp 1593098107
transform -1 0 1864 0 -1 210
box -4 -6 20 206
use FILL  SFILL18640x100
timestamp 1593098107
transform -1 0 1880 0 -1 210
box -4 -6 20 206
use FILL  SFILL18800x100
timestamp 1593098107
transform -1 0 1896 0 -1 210
box -4 -6 20 206
use FILL  SFILL18960x100
timestamp 1593098107
transform -1 0 1912 0 -1 210
box -4 -6 20 206
use OAI21X1  _196_
timestamp 1593098107
transform -1 0 1976 0 -1 210
box -4 -6 68 206
use AOI21X1  _195_
timestamp 1593098107
transform -1 0 2040 0 -1 210
box -4 -6 68 206
use BUFX2  _251_
timestamp 1593098107
transform 1 0 2040 0 -1 210
box -4 -6 52 206
use OAI21X1  _206_
timestamp 1593098107
transform 1 0 2088 0 -1 210
box -4 -6 68 206
use OAI21X1  _199_
timestamp 1593098107
transform 1 0 2152 0 -1 210
box -4 -6 68 206
use NOR2X1  _200_
timestamp 1593098107
transform 1 0 2216 0 -1 210
box -4 -6 52 206
use NAND3X1  _202_
timestamp 1593098107
transform -1 0 2328 0 -1 210
box -4 -6 68 206
use NAND2X1  _201_
timestamp 1593098107
transform -1 0 2376 0 -1 210
box -4 -6 52 206
use AOI21X1  _208_
timestamp 1593098107
transform 1 0 2376 0 -1 210
box -4 -6 68 206
use INVX1  _207_
timestamp 1593098107
transform -1 0 2472 0 -1 210
box -4 -6 36 206
use BUFX2  _249_
timestamp 1593098107
transform 1 0 2472 0 -1 210
box -4 -6 52 206
use FILL  FILL23920x100
timestamp 1593098107
transform -1 0 2536 0 -1 210
box -4 -6 20 206
use FILL  FILL24080x100
timestamp 1593098107
transform -1 0 2552 0 -1 210
box -4 -6 20 206
<< labels >>
flabel metal4 s 1856 -10 1920 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 640 -10 704 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal3 s 2589 1597 2595 1603 3 FreeSans 24 0 0 0 N[8]
port 2 nsew
flabel metal3 s 2589 1697 2595 1703 3 FreeSans 24 0 0 0 N[7]
port 3 nsew
flabel metal3 s 2589 297 2595 303 3 FreeSans 24 0 0 0 N[6]
port 4 nsew
flabel metal3 s 2589 257 2595 263 3 FreeSans 24 0 0 0 N[5]
port 5 nsew
flabel metal2 s 2205 -23 2211 -17 7 FreeSans 24 270 0 0 N[4]
port 6 nsew
flabel metal2 s 2013 -23 2019 -17 7 FreeSans 24 270 0 0 N[3]
port 7 nsew
flabel metal3 s 2589 537 2595 543 3 FreeSans 24 0 0 0 N[2]
port 8 nsew
flabel metal3 s 2589 597 2595 603 3 FreeSans 24 0 0 0 N[1]
port 9 nsew
flabel metal3 s -35 277 -29 283 7 FreeSans 24 0 0 0 N[0]
port 10 nsew
flabel metal3 s -35 557 -29 563 7 FreeSans 24 0 0 0 clock
port 11 nsew
flabel metal2 s 2045 1857 2051 1863 3 FreeSans 24 90 0 0 counter[7]
port 12 nsew
flabel metal3 s 2589 1537 2595 1543 3 FreeSans 24 0 0 0 counter[6]
port 13 nsew
flabel metal3 s 2589 897 2595 903 3 FreeSans 24 0 0 0 counter[5]
port 14 nsew
flabel metal3 s 2589 697 2595 703 3 FreeSans 24 0 0 0 counter[4]
port 15 nsew
flabel metal2 s 2061 -23 2067 -17 7 FreeSans 24 270 0 0 counter[3]
port 16 nsew
flabel metal3 s 2589 497 2595 503 3 FreeSans 24 0 0 0 counter[2]
port 17 nsew
flabel metal3 s 2589 97 2595 103 3 FreeSans 24 0 0 0 counter[1]
port 18 nsew
flabel metal3 s 2589 1497 2595 1503 3 FreeSans 24 0 0 0 counter[0]
port 19 nsew
flabel metal2 s 1549 1857 1555 1863 3 FreeSans 24 90 0 0 done
port 20 nsew
flabel metal3 s -35 1697 -29 1703 7 FreeSans 24 0 0 0 dp[8]
port 21 nsew
flabel metal3 s -35 937 -29 943 7 FreeSans 24 0 0 0 dp[7]
port 22 nsew
flabel metal3 s -35 1337 -29 1343 7 FreeSans 24 0 0 0 dp[6]
port 23 nsew
flabel metal3 s -35 497 -29 503 7 FreeSans 24 0 0 0 dp[5]
port 24 nsew
flabel metal2 s 381 -23 387 -17 7 FreeSans 24 270 0 0 dp[4]
port 25 nsew
flabel metal2 s 845 -23 851 -17 7 FreeSans 24 270 0 0 dp[3]
port 26 nsew
flabel metal2 s 765 1857 771 1863 3 FreeSans 24 90 0 0 dp[2]
port 27 nsew
flabel metal2 s 557 1857 563 1863 3 FreeSans 24 90 0 0 dp[1]
port 28 nsew
flabel metal3 s -35 317 -29 323 7 FreeSans 24 0 0 0 dp[0]
port 29 nsew
flabel metal2 s 1133 1857 1139 1863 3 FreeSans 24 90 0 0 reset
port 30 nsew
flabel metal2 s 733 1857 739 1863 3 FreeSans 24 90 0 0 sr[7]
port 31 nsew
flabel metal2 s 605 1857 611 1863 3 FreeSans 24 90 0 0 sr[6]
port 32 nsew
flabel metal3 s -35 1297 -29 1303 7 FreeSans 24 0 0 0 sr[5]
port 33 nsew
flabel metal3 s -35 897 -29 903 7 FreeSans 24 0 0 0 sr[4]
port 34 nsew
flabel metal2 s 893 -23 899 -17 7 FreeSans 24 270 0 0 sr[3]
port 35 nsew
flabel metal2 s 941 -23 947 -17 7 FreeSans 24 270 0 0 sr[2]
port 36 nsew
flabel metal2 s 1069 1857 1075 1863 3 FreeSans 24 90 0 0 sr[1]
port 37 nsew
flabel metal2 s 381 1857 387 1863 3 FreeSans 24 90 0 0 sr[0]
port 38 nsew
flabel metal2 s 1133 -23 1139 -17 7 FreeSans 24 270 0 0 start
port 39 nsew
<< end >>
