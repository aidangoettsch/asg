VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO basic
   CLASS BLOCK ;
   FOREIGN basic ;
   ORIGIN 3.6000 2.3000 ;
   SIZE 16.8000 BY 23.9000 ;
   PIN a
      PORT
         LAYER metal1 ;
	    RECT -3.6000 16.3000 -2.8000 16.4000 ;
	    RECT 1.2000 16.3000 2.0000 17.2000 ;
	    RECT -3.6000 15.7000 2.0000 16.3000 ;
	    RECT -3.6000 15.6000 -2.8000 15.7000 ;
	    RECT 1.2000 15.6000 2.0000 15.7000 ;
         LAYER metal2 ;
	    RECT -3.6000 15.6000 -2.8000 16.4000 ;
	    RECT -3.5000 6.4000 -2.9000 15.6000 ;
	    RECT -3.6000 5.6000 -2.8000 6.4000 ;
         LAYER metal3 ;
	    RECT -3.6000 5.6000 -2.8000 6.4000 ;
      END
   END a
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 0.4000 20.4000 9.2000 21.6000 ;
	    RECT 1.2000 17.8000 2.0000 20.4000 ;
	    RECT 6.0000 15.8000 6.8000 20.4000 ;
         LAYER metal2 ;
	    RECT 6.0000 15.6000 6.8000 16.6000 ;
         LAYER metal3 ;
	    RECT 6.0000 16.3000 6.8000 16.4000 ;
	    RECT 6.0000 15.7000 13.1000 16.3000 ;
	    RECT 6.0000 15.6000 6.8000 15.7000 ;
      END
   END gnd
   PIN o
      PORT
         LAYER metal1 ;
	    RECT 7.6000 14.3000 8.4000 19.8000 ;
	    RECT 12.4000 14.3000 13.2000 14.4000 ;
	    RECT 7.6000 13.7000 13.2000 14.3000 ;
	    RECT 7.6000 12.4000 8.4000 13.7000 ;
	    RECT 12.4000 13.6000 13.2000 13.7000 ;
	    RECT 7.8000 10.2000 8.4000 12.4000 ;
	    RECT 7.6000 2.2000 8.4000 10.2000 ;
         LAYER metal2 ;
	    RECT 12.4000 13.6000 13.2000 14.4000 ;
	    RECT 12.5000 12.4000 13.1000 13.6000 ;
	    RECT 12.4000 11.6000 13.2000 12.4000 ;
         LAYER metal3 ;
	    RECT 12.4000 11.6000 13.2000 12.4000 ;
      END
   END o
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 1.2000 1.6000 2.0000 6.2000 ;
	    RECT 6.0000 1.6000 6.8000 9.0000 ;
	    RECT 0.4000 0.4000 9.2000 1.6000 ;
         LAYER metal2 ;
	    RECT 6.0000 2.3000 6.8000 2.4000 ;
	    RECT 4.5000 1.7000 6.8000 2.3000 ;
	    RECT 4.5000 -2.3000 5.1000 1.7000 ;
	    RECT 6.0000 1.6000 6.8000 1.7000 ;
      END
   END vdd
   OBS
         LAYER metal1 ;
	    RECT 2.8000 12.3000 3.6000 19.8000 ;
	    RECT 4.4000 15.2000 5.2000 19.8000 ;
	    RECT 4.4000 14.6000 6.6000 15.2000 ;
	    RECT 4.4000 12.3000 5.2000 13.2000 ;
	    RECT 2.8000 11.7000 5.2000 12.3000 ;
	    RECT 2.8000 2.2000 3.6000 11.7000 ;
	    RECT 4.4000 11.6000 5.2000 11.7000 ;
	    RECT 6.0000 11.6000 6.6000 14.6000 ;
	    RECT 6.0000 10.8000 7.2000 11.6000 ;
	    RECT 6.0000 10.2000 6.6000 10.8000 ;
	    RECT 4.4000 9.6000 6.6000 10.2000 ;
	    RECT 4.4000 2.2000 5.2000 9.6000 ;
   END
END basic
